PK   �cU9_���P  �[    cirkitFile.json�}[�%7r�_1j_;�2���e�֞���� 	y�ӥ���<+�_2ϥ�$�ddEP��[]I~�����^~x��c�|������_�>?|������S�����Ï��O/O�?=�?���������_~���y����9i0tJ5S?�F��?�[ӈ�Cg�q��I���7�~���@F' s�"��$s�"��"s�"��&s�"��!s�"��%s�"�SK�@E��́� N�́��}�Q�!<WI��@w�dς�.���a�!<��$Cxt�I��,�n��Y�'³��N2���输�Y�}'³`4�S�}'³��N2�gA��dς�;���w�!<��$Cxt�I��9!�w�!<��$Cxt�I��,�t��Tt�I��,输�Y�}'³��N2�gA��dς�;��龓�Y�}'³��N2�gA��dςa���;5�w�!<��$Cxt�I��,输�Y�}'B��w�!<��$Cxt�I��,输�Y�}'³`�"��NC��dς�;���w�!<��$C����N2�gA��dς�;#��~������z���ǧO����_|�/��`�cc�y�� Fa�&�Y� l̨6��֚����Eivce���I��N�ڎ��'��Vǧ?���y��r�:���Y�`�FO�jz7�f��leg'7�'A�T��<�D�Dd68�Ӽj׼jge��|��Q�\Zg�PM���0�Ƶ]�(X���;Q��vIT{d68���j��jge��ĩ�]�k;Vv�K}PnS;�j[�h����R]ggk�!wd��;^�G��m'��'�kv�kvVv��.�QeN?�D��0��f~au-����7��9���s8^~��/�hf�k�����_X��l?權�0��ș�J�a��-c��>@Ѣ��k��d�v�sʑx_�F4s��)/?`��3ۏ9M�����vLB��T��0�J��᱘�9�朇�$���&�Ew}�4j��X4�ӲiaMR�V��&�&ɜ0���m*j���ja7��s-^~��/�#b��|��s�%�s-ɜk��f~a����s-^~��/�:c�*���q��vhİ��l�N5s�:i}/u��_�F4s�%�\&e����br}3H���q��ΝF�^[��t�3�i�MŜ�I�4��0�;#���2I�J���מaQ�VJ7�������<�y�t�Ӵ�Ո�bN�$s����������S;� _���Ĭ��������R�Y��I�J#�y��Ո�bεs������}����r��`���J�e�C�[75�֭�.�('ܰ��.�A�Ո�B�lD}�䕍�^�j|x,�g��s����������cM���0������<%��������ǜk��f~�$f�1�k���TWR����Ffit�ۦW��L�3Ɖց�.f�G0�5��zk:�1��F;����6N�h��@�G�_��V�²�5[��25V��q��᱘�9���/?`�NGa��l/?`��ua�s������i��ǽ�{CX�/���M���H6Z	��A3e�Ό�0)r����4͜����m*j���j��!f�3gx����_85��~�/?`��{b�s�����������<%�����3�x�g��^~��/��l?欇�0��1ۏ9�����l��c�zx�A�_*tk�N�H'�:�8�C�,���:��aN�s��{���Q;鉶���M�Z�8����l�����F�lg�EM�Tܧh0'L&JH�m*��aε�W��c1=s�e�s-^~��/��l?�\��0�'[2ۏ9���������̹/?`�Ne�s����R]�4+@�f��Ӯ�^���D'��9ֵQ����q��6fP�����ގ����Nv-�}�R��K�,8.�#�pvA55p���Y��׷��F���d�if9���ڡ�ut�����3{V��{�����շG���=��`��a��oO�>X}{�����s��ʆ*;��A��'*/���h}����/��'�/�m�h}����֧�=������'�/���h}���{���'�/�k�h�E�_t����Ԏ����6������n`;Z����ֳ�����n;Z����v�����Q�]XG���?u�>QѝOGCg���{���'�/���h}j�A�_t���y�i�V
_A���������V�2��w;Y'�z��Q�󍏪�o{T�|ӣ��[U=����vϻT����Ɇ*;��v�N\}��v�N\}��v�N\}��v�N\}��v�N\}��#�o'���'�o'���'�o'���'�o'��u\D��d���Ԏ�����W�����W�����W�����W�����W�����u�����u�����u�Bg��v�N\}��v�N\}j�A��N։�O�_t����y�95����]�͠�~������u�0���zQ���CUϋU=�=T���P���CU�U=�;T���PՉ���zq�����zq�����zq�����zq�����zq�����zq��~�����W�����W�����W������q������S;^��v�^\}��v�^\}��v�^\}��v�^\}��v�^\}j�G��N֋�O��N֋�O��N֋�����zq�����zq���G^�SS߮��J��%�>�I�4��n��'l�Ь�r?�;r�h���
�
2����q�_�f�1�J޷���]�,p�!Fʎ���ַ�-����^{D5�R�v����툪��#�z��@U�w����U=� o��ih{c�J^��y o�$�`>&�6D7�G%�&�K�(o߿G�D*���T$�ﴙ_v�w���7������Ah�6`V]ggkUYpj1́bBm��A1!����P�sh���Zs�c���8�z�3GU�w����U=ߙ���P��#������1$�~����'
og�	��WP���'��RLs����*�JP]�`o�O��M�Bu����	Tv��0�I吓�W�<9�_�N��|�ܻ�4C�f�s��M#}� %r���BU�7�:y� �%��E9��B��V}g5���b,Lu��L�3DF̄_��_FfN�_n3����"׿�~���2�$l�/��/�N�#�2��d0D����4����4-~���p!����>��;�=Q�w�{����D@�ז���eg�2��"��{{��3>���savʍpU0�u槑ӭ�����ri����o�s���_����E{�I�����B����n��b�̛#���%�ۓx	T�y����4d Ch��������gB�Bm��-4*�P��-嗩���@����T�Ζ��"7��i�?�=PL�q3j�A�R,��3͞� G�e¼p��Y۪eoTS}'P�T�U�T�	�1�w"~L���S}'n�T�	�1�wvwa���(�PeG������D��%���D��%���D��.��O��^���O�{D��.��O������D��.��O�����������%P��/Q{�K����w��>Q{�K����w��>Q{�K��S#?����@�'�o�p	T}����@��D��.��O�������ԃ����%P����;\U��?Kԟ%���g���D��U]N/O�������7?��s?O����M��������. 7x1�0^�È	H�!FL@"���0ba����cO<���D��a�$�#& �x1�u��E�ym>��淁�qs!�u����6�ͅ$ֱV&Nl��8�XǄ�8��p`s�\Hb�f����%��B�;'���/ g��͏s!�u~����l~�I�� L����d��\Hb��a����%��B�S:�����B��'����6?���8�X���8��q��ǹ��:G�ĉ͏+6?΅$ֹT&Nl~\��q.$���2qb��͏s!�un��ߘ8ߠ8��l~�I���L����f��\Hb]?�ĉ͏k6?΅$�uLS?l~ܰ�q.$���`������B�&N|��|ӛl~ܰ�q.$���a������B��&Nl~ܲ�q.$��Ab����-��!�+�9�ȣ��w��a�ʵ54T���p'��r�$��-P�+T�*N��]e���
U�FZ1�U��\9��J����W]E�5�B��nc&��*z��r�5ŕn[E���^kp�*\��Ӓ��V�k��y�LqVWŮ]��\9��\��U���b�\�
װ&�Nb��bb�l�۰���m+e]�Ү:y�I��N�U�-�a֚ױm��갅:lÚ�:����Uau��_s�i�:YX��f�`�:���Ī��:l�^�:����Uau��w�1�@��,���Ӷu����Z\F���%����WzqM,���l9���{��ضN^V�-�a�\ձm��JSbu�2Y'/�u�*l�۰��m��eU�B��w~rڶN^V�-��2�N^����˶u�$[#���d���
[�����{Nۦ2���˒l�P'/�u�*l���{�m���keR���$[#���T���
[��6졮c�T�à�:yY�-�*-V���%�r�rڶN^���eU�B�ao~���t�[��6�1PǶu�˪��:l�Y	ul['/���wwGqڶ�|Y��ZLs:�+¸l[c*�ЌiN'ɖn���L1��3_�`��i�:y����Uau؆3Q�ض�|Y�P�m8ۥ�m��eU�B����ON�V�IVi+Y�-=N�^��e�:yY�-G�P�m83��m��eU�B���:����Uau؆3��ضN^V�-�a΢�c�:�eU�B��L�*�5u�*l��p6X���˪��:l�gul['/���g�ձm���
[H����N^f��e	��C���:��t�G�c>��e&�tXP���%�r�rڶN^f��eU�B��L�:����Uau؆�%�ضN^V�-�a�Ȭb[['/���g}ֱm���
[H��Ƿ6�t8�[gc��f��}�$�,�r�a,���㤚�
��r[=�C?��=�Q2g�Dɜ&{%s��A����Q2geDɜn}%s�A��	�Q2g>U�xyԛ���(�~sW���Qp�ӣ0<�]z�GŹ�8��0�`�n�<
ã��]�GaxT��q�(��s��uyT��=�(S(���ܵzGaxT����(��sW���Qq�"��0<*�]wv�)"�Qq���0<*�ݶu�GŹ;��f<*��u�GŹ����0%v<*�]\t��b�J��i5x�]�΍h,��{W@�U�B)��R�
�(JQ1(��`P(<z):=J���T�$^���p0<�-��`x\���h�<���Qqy, ��yT\���<���Qqy, ã��X ���Qqy, �J�<���Qqy, ã��X �G�� ���c8���G�� ���c8��pY���c8��p0L����c8�
>
ST�S��[_Y��5���'�k�Z7���
��aJQ�(���Q(E�P��E��B)��R/
�G��	�z�#8��G&p0<
.�L�`x4\����<2��a��<*.�L�`xT\����<2���Qqyd���<2��a
%xT\����<2���Qqydã����G��	SḌ����G��	���#���G��	���#8�Į��e�s+}�e�C�[75�O���rq��5���8�����I�Ce������h��+�5F'�y��e.(��f�i05
1��$����8�Bӹa�U]���AY�ؾ�vL����A̪�وFfn|�o]��d�t��%�dr��-�P��
E����8��m�9��h�-M�����{)�u��-(��]P(E��P��Rt0(��A�;�Eخw��t3xg'���;��n2B��9��_ 
���(�bK�P�_@ߎ�<�C#���l�N5s�:iu�Cg�^
�R��_�_�����uZ6-L�s)L��\P(Pji��F��T;g���+w�c��a�Ah�b�U�����.
��F(����� 8������~�8��`}a���m5M���ž�R��P(E��B)zLJ�c�P��R�*P(Ť�R�)p�+v�8������ȷ<�>��
���d�?�i��)l�h':��t�T�{ �=
E�foMgA4������a\�$�VK�� eO�B)z*J9}Ġ�-�f!�L�4yΓ�>��S�'C�n6�й���yr�X�
���P�vA�#!Jy���aZlc��(|��m3M!/�>@�{�*yJy=����R^M�Aᱮ)�0([��P(k���TO@��fQ����o��eIQ]���@�O�`�� �G��U�(��j Ly5
��ӕ�LyM���`�*y�,��`�}\vL�Kì8���A�R`xT\��tk�N�H}��| �lͲt�[@�sϽ�CQ(��Rt}`;7u>��f�Eh��;h��ԙq�ۺ�|߂B)�
��F�k�MK#�4��mӫi�M�|�#Z��F{}.
��F��ɥuV
մ�y,Ƈ�m�7
�E<�y���ޗ�B)�
����R,>\n�4{�A�>�6a�2`tֶjAD����Š�#`J9����J9~���/�=`P�K�1(���:&���Oã_D���Q0"F��h�OãbD��a��<*F�E���Oãb�>Q���DQ�.���DQ0L����DQ0<*F�E���Oãb�>Q���DQ0L1���DQ0<*F�E���O�u��Oãb�>QSbǣb�>Q���DQ0<*�<*�<*�<*�<*�<*�oU�����t��ҿ�����;<��4<���4��x��/������XǨX1�u����X��X1�u���X��X1�u|���X�Y1�uܒ��X�@Y1��x*�����|n��o���B�acNl�؜7�8h�pb��������y����6'΅$Γ <����d��\H�<=�É/������d��\H�<�É͏K6?΅$��C<����d��\H�<s�É͏K6?΅$�sj<�8�Wl~�I�g�x8�����q��ǹ��yR���Wl~�I��[y8��q��ǹ��y"����l~�I���y8��q��ǹ��y�ߘ8ߠ8��l~�I���pb��͏s!���Nl~\��q.$q^W�3������B�<����a��\H�����&��&�7l~�I����pb��͏s!��b Nl~ܲ�q.$q^��É͏[6?�C�����y�?���~|��??���W�R���'T���p��]��]kp�*\�IV���b�\�
WqRU쪪صW����]U쪫صW����AU�j�صW����(U�j�صW��U��*vm�صW��U��*v�صW��U�\��*v���pk��$u2�*l�۰���m+e]�Ү:y�I��N�U�-�a֚ױm��
[��6���c�:X�P�mX�_Ƕu��*l�۰���m�dbU�B�a/F���ƪ��:lÞ�:����Uau؆�1ul['+���{|�L,��˪��:l�^�:����Uau؆=Wul[iF�ҔX��L���d���
[��6쁫c�:yY�P�m��WǶu�*l�۰'��m��eU�B�aoe���˪��:l��:����Uau؆��ul['/���{v�,L���Uau؆��ul['/���{��ضN^V�-�a��ױm�Պ��+���T��L��˪��:l���:����Uau؆3�ضN^V�-�a�J�c�:yY�P�m8�m��eU�B���:����Uau؆38��V��˪��:l�Y"ul['/���g�Աm���
[��6��RǶu�*l��pFM�V�IVi+Y��L���t���
[��6�TǶu�*l��p�Q���˪��:l�Nul['/���gQձm���
[��6��UŶ�N^V�-�a��c�:yY�P�m8㬎m��eU�B�ᬶ:����Uau؆3��ضN^V�-�a�Ϋc�J�|T:�N^f��e�N^V�-�a�2�c�:yY�P�m8���m��eU�B��l�:����Uau؆32�����˪��:l�Y�ul['/���g�ֱm���
[��}�+�,�r�a,���㤚�
��r[=�C?��=�Q2g�Dɜ&{%s��A����Q2geDɜn}%s�A��	�Q2g>U�xyԛ���(�~sW���Qp�ӣ0<�]z�GŹ�8��0�`�n�<
ã��]�GaxT��q�(��s��uyT��=�(S(���ܵzGaxT����(��sW���Qq�"��0<*�]wv�)"�Qq���0<*�ݶu�GŹ;��f<*��u�GŹ����0%v<*�]\t��b�J��i5x�]�΍h,��{W@�U�B)��R�
�(JQ1(��`P(<z):=J���T�$^���p0<�-��`x\���h�<���Qqy, ��yT\���<���Qqy, ã��X ���Qqy, �J�<���Qqy, ã��X �G�� ���c8���G�� ���c8��pY���c8��p0L����c8�
>
ST�S��[_Y��5���'�k�Z7���
��aJQ�(���Q(E�P��E��B)��R/
�G��	�z�#8��G&p0<
.�L�`x4\����<2��a��<*.�L�`xT\����<2���Qqyd���<2��a
%xT\����<2���Qqydã����G��	SḌ����G��	���#���G��	���#8�Į��e�s+}�e�C�[75�O���rq�K9�F��i������h��+�5F'�y��e.(�25
1��$����8�Bӹa�U]���A)rM߃�U������޺V��,z�d�
��K�SB��$e�ILm��)�F�ni�������Ki���oA��B)���c���A��
��I.�v�[Ʀ��;;�M���ht��-�)��%J��Q(ŖF�[�o�eڡ��z�qK���o����3e��P�v���K�}^@qиN˦��� �i_#
��K���r�1������*�Yu����P�1��F�0��[��}�留3M���8��vQӄ��0(����F���R��(���D�=&
��U�P�I
��S�T�$^����q0E�N���i&�w��x��}ډN*1!<
�hJ����tDc@��ى���5N�h���\ �R���7*��7�<9�(;5z�1t�f�����'7���Ơ�[�R�
��.���n�i���o��a�v��4��D� mFd}(��z
Jy9�����c��Z
Jy)����R^H�A)�B��I�<�E��G����Jã`�*y����Q0<*F��G�0�`#Vɣ`xT�X%���Qqy.zЭ;A#a���򁴳=4�ҙnq ���=7
��JQ4`;7u>��f�Eh��;h��ԙq&ĺ8J�P(�7����҈�,��{��j�}S;��ց@�
��F��ɥuV
մ�y,Ƈ�m�7
�E<�yA�
��F(����X|�ܘi�(�}Dm�0e��mb>�R���7*�^J��bPʞ�Rv��r�A)�r�R�xyԋ��Q0<�ED�(#"`��0
�Gň��yT���Q0<*FD�(#���`xT��'��uyT��'��a
%xT��'���Q1b�(
�Gň}�(#���`xT��'��a��yT��'���Q1b�(
�Gň}����Gň}�(#���`�;#���`xT��'���Q��Q��Q��Q��Q��Q�}��~����/�������q�χo ><���<9����������<���|�-er�e���� p�|\�1�$.]E�����@�[,>f��\�v�����)k�@Y9�B���^�B�h��uo*�i���*D�l/��Q�M���(��
n��F�CY���-@��
r;��AY�p��@r�K:H��@p��
r�9�
N*���$&-�&��T$�*�2
r�
.ZA.�%QѸ��j�f���\nK���p�d��������d{�&�
Q)ۋO3T��8hTPFA.�bB�`�!�����A.�%��"��ȝ��v�t��!���UԔȜ��-)Γ�_��`���&����uC��1�q$*��!O�Q���wi�1�AH?�H@�i��i�lZ�o���c����c�N��)5���'�t�>СQ�{_)��L��[+q�
$(��&�	���6�2U@g�=c���W�8�3�?�e��L#�q�&�3�5&茸�v�*StF�3��~�	:#�y�]F�����,�.�_e2�Έ{Nb��~��	:#���x�W���b���%��L[�q�^�2�5&1脘�2��7uJ��{�3C�	:�<=�!Nw�s�=�$N~�C9��~J�kL��w(�ƌ�>�_cb��j��z+Q�I�B�-�e��L��i��y������������iY�?wzy:}}�����Ǉ繟�'_=��Oo�� :�X�� � C���"2�X�� � C���"2�X�!� C���"2�X�8!� C���"2�X�X!� C��-T���=9�'��J��Sf�<|(08Q:�8�sC���G����1���*_
Δ�!�g�Py0�S��O��|��G<��2�S��O��|`��?����!�G6Qy0�S��O��|h��?����!��VQSI��)C�΢����9R|��)C�����`����1���1*��)C��?��`����1<J��#ܨ<��f�tq>D�ʃ��jJ��c�<��f�tq>H�ʃ��jJ��������0�S:�8&H���O�?�c��q�T�P�P��0�S:�8��H���O�?�c��T��2�S:�8�JI���O-�?�1��	�y��#�ݬQ��I�����������	��m	[�$<`����I2�O2ۏ�0��"l�-�߾��z$�ۏ���%ZW3�S3���0��8D�l�Iu�4kD�֍��k��i��������Y��2ۏ�_�!s�� �s��dsv���m^�䌀��89fs:fs��f~a�$wh��X��!p3+?�mȞ߰'8�p�8���03n�a�-�y3�f��janrg3������(<6,�0@L��	C�0��Yp�1���aXp�mC�T��!p3��a��D�Hp�31aF@�r�0�C��̝��7*24l¢��s'51ÍH�7��ۤ�93C�fv�pې}�}"�;Ǒ�9���q�7ð��ۆ�93C�fx\�9�&��3�a��s��Q/[�*ҹ��M���Ny$w�����a�c�(��Ȓ8!�L���Ny$w�������b��)�QJ�h`&	�Tp�8�;�af��a�Al�%qB��0$S-PX�F��Cqg@1aF@�rg@�;bf��~an�&�������6��af��>mnr�8�������ǆ��8��+N�^��@~�&M$�-4�A�]�����s(���u��3�p��h5w������m�=������$�mȝ�03n���3���aߘ1��iKD���Mʝ��7 Ny0��p��;bf���*�6�΀�7�p*��3 f���0�h�mC�if���0���lCÝ�03n��$!nrg1���a8�ۆ�Y3C�f(�nc�!w��0��:�?��g�Wn�Mʝ��7 �W2���Ǥ�H����0$S-��Vw���;�afN;�V)w������ڸmȝ�03n��9nr�8���a8!�ن�;�af���~�6��q�B��&�"��QB��'�'��J6A��-�'�)���5��u�f�`���'��V�f�����Y��U��Ly�~t�����ɺ�G'���d{�~t����ɱ�G'����zT?dR_�w����Z�� T����0���( U��eiGȾ����^�� T%�7y�*1�;�( U��mUG�4�������e�㫔�P�_^t������� T%���*1��( 9B�*1�=�( U��}-G�J�oH9gS��Ir������ �d����� ;J�`���V�������V�2��w{�*���
P�wD����T�	���( UG �����qD��;~�� �
��Wq T��8 �
��U U�{�*��Ľ|@��T%��8 ���U U�{�*��Ľ|קQ����� ��2U�{�*��Ľ|@U�^���*q/_�P����� �"U�{�*��Ľ|@U�^�����J��Wq T%��8 r�BU�^���*1�R�(�������jҍ��f�M?Y�X��кq@�ę�;:D�ߑ!���
Q�wD����AT�	���(UG���T��e�8 ��2f U�{3��½�@��^ƌ�*q/c��}!U�{3��Ľ�@U�^ƌ�*q/c��iT%�e�8 r�LU�^ƌ�*q/c�P���1� �J�˘q T%�e�8 r�HU�^ƌ�*q/c�P���1��l��2f U�{3����(q���J_cY����M����Fv �\�pòf��˕�O�<1�K��R�~�7â|F����5F'�y��)v-.f�EN�BL�o	}�{�4δ�tnzmUק�u�;HÍ��A̪�وFfn�R�o
��d�t2�2�Pp;��η������(K�qS�z늱Ѳ[���u3�V�4��G��1���9P�w<����A���;��;�"l׻el��������XF7���r)uK�Ns���4'�~B�*׷�2�Јai�{۸�S�ܷNZ��Й�ut�:(��q����.�wиN˦��� �iu��.v���6��������z�:c���Ah�q�U�����=d�,\�e34
.񲙦��A���|o�iz�>1��ζ�����ʌ�Pp��J
���U�ɢ��8YT�'����dQ�w�T��U'���i����x> U�{C��,���L3ɰ�����M>��;�NtR�)�T&�E��_��|�(�����zk:�1�}�����'A�Z�l�T� 3/��K��LD���K71�� AfB�ɛw���1��=�غw�i���ևՓ�Ɣ�2A
n�SA�߱�~�:�
�7�ݍ�0-�1��>�ގ�����H�����eL��� ��{�0��`�S�gЁ

΢�<\�eĆ��b�̧��s1\�oᤈ�Cpx	��qd8�D/Bz_��wL� �  �  �  bM�h�Vh�"�#ﮟF�:͍����./7������[^��ef�G��L�[v�F���qg{h��3�� Zץ��L���t&�G�%�`f�l�\��N�f��(;uf��I�^6�)��/�
.���>���Ffit�ۦW���|�%Z"ٲ����|�(��e!�;���J��v9�����F����0�yI�l�D�%��Qp��ʌ�u/�����L����CzFZXgm���@S��c����{���^,����`��9mL��@SoA.��^܁�Y�T�� DP5�� �*��Q T�� DP��� Ⱦ�����( �ww� �J��A��*qw!�O�*qw!
��-S����@U��B U��;Q T%�� DP����@��J��A��*qw!
������8�����( �ww� ��
U��;Q T%�� DP�h�J�T%Z�-U���D{V�_?<�V|�N/O'���ᛟ0(=|��C8
�=a�-�I�y�0�X��H�	C_��:.�.�[�����V몡u%Һt]<�N��S����:_���YWݬ�8���::�NѬ�>��:����i��ܺtx]��.�]���u�{]���75t��Cj�PC�&�0��	5L�a֗5L��?��jy?���3��?���ޔ���3�)��0k�_��+`���W@����YL����`�e��A,vM�:f��{b�v��R�9b�dT	�N��m�����_�j(im�
��+�6�^��ƈ�z�yK��t�g�u�7��}��/�jת�]�a�v���꼹}q��M��P3}�[�?�*f*.j)̔V\	15U�L�D�0�o���%���I�%Bj�PÆ6�����>�z�?�/!<�տ��\�Y�b�7A+����� �#݄�ӓw����[�b�d��X\d��3�\8L"WnwCaG�h�;rbv6��N��n{7b̮��#�n{we̮˰C.;!�����svD�i]��5r��r�A��C.����J��v���~�����"�3%���
�?R��R�������\�v���_�Į(�\W��I"ז,��)��I߄R%��z
��w�Rt's=r���.}�2�S �q�lW�be��@�â�+�.�Q wUq�K[.�O w��m�_����	�ff�R+s�r�.�]�t�~���\�r�~�����:f����BI�"6�6�C�[���"��e6 �z�drn�����%���:r���ɴ	2�p����&��6���1	29'�<������rU�K#O�"���\��4�t.;[b�s�ȃ�H��"6:綑��v!�lrnyi�e�&緑g)�t�F^'�^��|9}��S���&��u~��`��#qy$�G��HƏ�告��#?2�G&~d/�l���<j�G��Q?r�G.z�W����f��Tp����A �\-�I�j�mW�@l�b���*��f��.�j�E^�"c�țNb�ȫ]dly����"�v��]��.2����E�v�W���.�j�E]�b���]Tlu����nPlu����vQ�]��.*����E�vQW���.�j�E_�c��]tl}�����O�N���O�S�<�?/O�O�_^���IO0v�N�Xxc��I�
=!����ɪ�<��篳���i^^֙y�C}�	F}���!���~xY�id2�̭7���KX�����?<?�8?�<��R�?��9��ЅxC~yy~�&k?��O?<�G��k��t�G��������O?���?xЇo��ӗ�?�2?������|�����>>���7/��o�?���.����y~�����^i���_��>���?���:�V�֏O__��A��	�	��J�����:o����}Շ�);�H��`�v�}�(ǡ1�9�Fe:1yN�������s���O��>��gF_���O�9�m�l?�^6���C��LV���G ?��6���?%�H��P@�uݪ&����Oi.��!~�F��_���K��?�"H'Ο��k�v-gΌZwf�\�'�_J���]-u.��~J	�������+��^�Ɯ�Y���:[©K1u{��I����ri�r}A�l�OҌ和�riFbeJD��'iF�rIFq�$#pg��nu�x�d�*�b�(�fԞ��6b?I3J�K2��e����|� ?��0*g�o��>�+��A�w\,I;*�f��o׹�+��I�O�\�P\.�H�ĥ0[�'��%�%��Ҍ`e.e�=&��%�%��Ҍę���}�*��I�Q�\�Q\.f������_�N�O�6?9G�>
SC>���"!�����)�}�m߆~��f�f��614���f{ƍ�Y�v b؆~��A��O�7���f���[��?�װ�Z��t�����>����"� 	 fS�e�i�*�C������(�$M).��(�&���w7N�4��\�Q\.MH���A�PT.C(.�&*j�sD�-(�\�&����3����u8�!K�O=I�OL�OL�os&M=I��fH%
�I٬�OҤ�R��iR:k�ē4��`�T�`���Z*�$M*.�!�(�&YK%��I%
B�T\0�>Q0�^dM�x�f�(�f̰O��W}�*�넋�C���>�3`�n��-�ҹ�����9-����A�� �� �����қ�?��'��{��EF��I��ص�З���'�a���
�:y���k ҝ;A�nO�}Ǩ���e ϧ�gC�\��O�^ŵ�>׸a�(���ߪ܆.�3������mso�)��B��[f��5|�H��2%ύ�y��H��ރ9�0��j�������w׿���R*J�u�.+)].!�t������(]⭊�%R"J<k(�,!�tA�rP���;�.�R�We��ګ��j���t�v&�u'K޻�t�;��.��^�)��.�p�q��A������F���0����O��_�=|�V�Z���(�l��c{7��ɩU0A3�fifP��l磙E�L����u�"��B���ս���[�Mb��6b0T���Ah@�G,Wȵs���h����d1`�
��:ٮ��2P��4�/��Bw�>��cw���
a�5�c�3/����Ǿk,�0tzr��[!���B�mw�������.$�ԃ_`����Mw���?{?�
�S�?Ȼ��A�MLӆ%nޣ�M+d��jt�,�����uB>�*e¨]�my_�~�����{^�.3�u��I��.�?�ӿ6`��~��������gv-j����,p�^���0	c��l�W�h}_6��;���t3ʶo���<G.u�B�ʽ�-}�K�������u�	n+�R%���B�5봾i�\J�>�prЪ߂�~	/��Au�>b>�O}��CV�5�m1�[�Mz�a���h�n]3*��jAM��g��Iu� Fb렄�AI*�AX#�8���(�����p���Q��(��Y�->���F��"��� g��r�F�l\�N��繑֊�}��N݉ u��V���l�U�� r��fn�͓u�j��ߔ��%��R���o5C��P�X��5��oM�]n����$t�^��k���G�>v�Qץ����>�7�]��+e[�Y��)�b���?��MB8P��sP,jVq����b������>A��y{r^$�u��<����r���yV�׵���Ī�>�k���>{��>��^w�Ȗ�>�b�3�D��Z�l�ρ�~9��ߔ�`Úds[�7��+��:П+������Z���t`x����p��x�绝����Rދ�@֓��9v�_#�#�|�?���톹�eۦ5�V�>��F�Pc�z^�R�m��^��[9�i���7巗D���߅/��\�(�F�h�aq��f��)�Q�*#L�.�R�1��߻�����]{~@7\k}��}Bu݀���UpO�����z�w�s�n�-����%f_7^\�:\�M��zW�-r�oc^�[������3bՁ|l�s���n�����f���?>==���|�����z��v�7ط?�����
������������N����_~����J��Џ���积��x�����~%�-����mY���¯��c?޿y�G��n?��a}����7����>������ߜD�=|�(�hY�7�����.���_���m������Ϗ}����_��c�?vm[�[��]���h��
�	͆=����aF,ш����S��>�?������o�/�1i>��H^u�=>R>\i��Zh!���b��1�.V��1����0���mlj���%�`�A�{��>AX�2�����K�6��K��ɹ�����z�zUs�����ۓ�"�[��Z�s*u��nO�K���K�������޼���n�V���p����沟C�ؾ�9�V�+��z(e�<o�	�R��ڼ�c����^�ϓT�mo�y��+}"/h�߿,���������o^�����'��.O��>y�0�?ŭx}���I���Xa�'��?��~m͓�ْ}�0ߥ��ɔQ��>��p�|������l�E͕7�-X{�p�p
u��P��V^M�1�����fcI�3b�Y:V��*w�F�\�Y�!�Àz�4�x�_B�k�wTm�Q���wxo�`����w%됁�SbiZ�4�@GC�K�p#�]xs߳���#'�u���w->v��z������_h��:���� ���!������p�wIn�R1S�X1���sz0��}a.�B�`�W�nG�nV��[�)xY��]Ŧs/���2�L9q=�c���H�������a(�r��5��$�.W�ȶ�.=�<��6֞+w����n��y�§S7W�.p9�L�'�"����%b�nKDM�-��@,�m�Hu��~�%�Oa[b����^���>��q�E��'g���V�c�MH��ȋ׹�́'�L�x�v�g���%L�.�h�t�����b�$�%��.K8].�1�&��t��M��?�t�����tq"���b�{���vI���.5\�X��d�XV�b�J��bէ�şQ���)�9��>����`a��-�Է�^��V�>]�[���B�#��Ga�t����0�c+��N���
��	�!U�}�]�mך�y�Q��n�D�k�s��Vm�y���`]�t���� �V�q1e>*���>���8���G�7��$��}��'�����O����s>�?��y=���Յ#L�s���ۺ�������<����?<�//�������#�/�П��A�������.�T���>|��������yZ����m�<%�ȗw����Od%���"��?����a����{G��~�Cx��5����ͷ����{2�m(J|Hk�xx-��ۿc�um���j�D������_�8�u��߭�9u�UәO��u���ٕ�a���Ɔ��:��M1�Pw�d�.'n[(�n�Q��e���:ݒ�X���0�����5tw�0������d�XZZ���z�q-i!:N�u���nt+�t�ֺB�*���"iE�zG��ԬRzw�x�+�vX����'�5`�)Nor��o�&�w���r6y���&7�����q���6��Ru|�����)�G��~�:���r�2�t��r5��{^	�wz�\9%��{XB��(����Jm[��B]�녴y�:��QB)�%�rAHQ��X�j^��;�����I�=(���y�t~	�����缽����seN��Q�(�rJ:�JU�:���:�{���s�O��Q���m1����V̽�Tσ9��$X��{��9��q�!E��x�}K�]r$mS
;��W�L�x�ۼ�W����	�������$���Bo�{S�I���{#d�3��K�ycyl��]\��ݣ�b3�.M���Ū�(#rvp�N_q�+c���m�M��k�m Y#�������78@���鑀Ѩ�{[�����!��ݾ��>@���l�6�A}��bU�n�y�̑�R���pe�Rt����S��H޷���׍2!o���-�xW�榯��?*9�ܛRU�s�iG�_�~ot~�+cs��]^#�XiuGύ1 g�&��_�u�x���6=2o1�w[?�����o�w��*g[ӿ��fl�̇}��U*�n�B� ���{P���{�[n��^��il\�*�s�)�/1���� WFM��^��:�b5| ʈ���y�x���N���o�M��Z��[�.�@��/0'zp���� UN��c���&�o���K�W�O�m�+��PLi��wB�����:�T����픜]ymJ�m�x-%�<�Tfw�V^H�%@�r�k/�9��Qf=����;:�}�PmK�=/��R�zZ���m�h�gZfn���2����%��(�̎pC�� �wn>����� ~?t�,֥]�����RQt�qU�{`��W�v#	n�}�z��ͤ�WN��q_,���td�b���i},�l��ԇC���[���[���/�k��v&d1�:|��(�Tj-?c����q�W�ӽ/�G�������P�X���$ȳ�j��Q�m�qi�}פ�ĭ��8m܎x��/�bXm,�S-6rE���˿Z��q��6�{����=�~ﾘ���vȷ9P��p��֜��%5��[�9�0Xm`�Ή�p2{��>��eZ�H��6�z��E0۹����,�Էnj�[
�rq����{�D;��sj�~$�f��L��R�1��W
=&whBJj�/�`3,�ǃJ7�����F'�y��ĽNI�w�����Iѥ-K�Hg[*��U��T��P@L�o	���zi�i���0�ڪ�疎}�t�\9���{T:�u��2�hQ�i�%��8��Q��C�h����w8���s7˝��-�Qյ�����,�1�W����co���.�]��Q���5f�r(3��!Y�n���'�Q�8P���}'��*\����ŁN��#&BYq�S�\��aܚW���G$};.����0H�qK�3ɾu�ꮇ�w���.`8��3"��`P��>��1��R�T[v��C�[��>����˿�/��c����7AM_�<��y��������?���_�?	/��_���PK   �cUs�7+5J  dK  /   images/6c71542d-16cb-4630-930f-71c4de5e1144.png4�4\�����G%�F���w� zｷ�e�D	QB�����+��=z������]ks������s�Q�*�xؔ� O^NJ��|��` �_Q3?� y)q���m>�Գ�LWm�5��G8�� ��0P�����h(_׎��hx���๓}��2�Y2���e�`e�e���Kw*�/��|b��G��,�\*k���-/X�F��fg��œr�z�cvvJFK�G/�/i�)m�b]��8�X
�LTjYx�*?>��98����O"2����.d+E]r���q��JW���5,�3E�G\w���_����� �Bĺ9���� !A���7�D�L�2`qx�^2b��z�-|�_�Q��o���O���|�w��o2r|u��؁�P,$,��~��v�7�5==�ʕ�����I���1�B'x��G��'�w��*��#N����G�vW�)�S�J�К�V�%�0�=^뽌�S�13�E�j�^Tj�i�xJ,_3��������T��ٞ�Rd#%*1]{<�+KSH�������`)\�}�^�X&.�.C�f"��#Dj@���a!�B��L ����ecŇ�X�\_@買Ox��-�C�����?����dʲ�J�qQ��s�JC�е9���tx,xXb60u	Ȳ�l�Lˢ�:�l
�Ð��ق��}ǿ��Yn�x�t�E^�M��x��-G���M��άG8�jε�:��C��#�,t�H�M�Q~O���Q�)��%#�!���2�cS�!)�����k�l&m��%�� X�)�t�琰X2�_�N��DE��W�������(�]����R��TI��F���Q��A	�
��)�)/L�<�٣�п��yR6��n)R���D'�-�G\
���FF�K�Ă@g0�/"��9�	�M�#'�9H�a�
B�X
w>KF�"	�|s��/iIġA���a>)5�:뿦���[:y"�B"����N���/$5vq!��}�Y$>��X�3�CF1�y��h9�T#���!� h��+����ގ\WggЙ^�E�-����]�ȂrO�Q�����#���:NSA�Q���|Y�,	�����Rj��[�W����vHpc�z/�4g<QZ�v����&�^�Vɭ���a#���(�|�D�<��MQ�KO�Ѝp�/ �l����Ѝ �d+��ྉG�O��Q��{��ڣ��u6\�@B@����0�g���㒒��QF��c��
MHBQO��3�V3�rP�� ����V��J$���fvf�����v�Y{�{~�Ű?�������E>�=d
�=hh����I���Ě��$�/����š�6�:k��D�0�U;��`�e��gV71"�qq���O�,�ظ������;َۖ�E#�3�=乚����ԭ9LZ?�˾nP�6��e=F@$���'�����`B1@���a��C��4	M(���g�1�Kq��t�-_��,����pV��7$��铂��u��)��eɌ����=���m�������II(8=33�Q~�˼F�~�/�g�K�PxPI��y�6n5[���i���X�O����ߑ'���'�à� �����3V �
��F$j�ö}&=�e(!��s��M���&8���(Rjal#Pi�4���O�>%�|�jm��7o�s۶|�-��w�}�7���aގ9��xh�r-�H�L����=<ʪ
@BD�j�C�r޾�5ȱNw�#[�S>Y�b�I��������V��[���|�b�����=_�kX�Á��FpI�����V-��-y��B����D����^L�4-�G*L����pz�1��
U{�^��6)#g_L��B��['�D�Li:�aAU��ɚ�I�I+@����ދ�4��ޑ�-��؎��M��L|A��"�É������ҧ��T���}*�#O֪�x���ٿZYZ�>�$�������~�<lc�w���]��TW�Z^N0�ZZ2�̇ȧ*�p����;Sc***:����hkk��^��?�%T[��;Ș�������k��g2*Q�����I�ʲ�I�H�(�D��mN����7���X�j����M������(���Qn4t��Q�����}���������@�?�̉������;��&�wڷ�����ɰ�I�m$���2*ʠ�:�Zh=�MX���e&���C��X7 �Kz�G���O#����６|���������m/?��l�"�
tIr���$=�е����_��m���C��^Ӷz6��+^���-G ���%�"O���_鱧%��ώ9��r�!����d�; I���|8˗�(���8���EF��׎W{>��Ńl2#֏{��^szdM�FD'1i��	j�V>�*)Y��yq1��8�	��?I�Qz�C$:��h?�􉅲�_vb/�� b?��m	8*�䍳-������@�{��z���ͪdԹ].��;{���X/V��_�*b8OP�(j������̱K�w܌t�Hjz�:�����Ҧ�5�m9���O��Z=,��X��\�����}�W)m�����CKPe�PS"�N��Jq?WgG�v��kt^E�} ̩����$�R�t_2��QRRv���!tZ[G'x�G���| � ����˥֝�ʳ/5���XP��R�/x(&�ݟ� ��xJͣٴ�[?n�|��ܪ������l�bZ���;o(�5tx�b�x3k��I�Q��U��c	GD'���!F"�Є ������}���8��BP����4f9e[w�o��@�l�&��E�1��p�˷�HQA�ֲP��S��P���n�"%R�Q��\ڐ	(��ۘy��3������Ue;�?�u��)�-p1w�s�Dh~�	���:��;J�VF,FR�}�B�.��Z�Q�g�9���O��!Mr5^Х*V�غq�}�g������d~�xA]����H��ː��w�Nf2 c����R��l����m��]���oyےV�:���i5��D9�1@IYy���X{��>ӹ*����D|��w��¾6}k]�5a߾PI>!�(��B�d�jg��/��P�U��\���l�!v-���1�~�{	C�����7�tp��ফ���T�|P��?�DL���QSS��8bBt嶫������~�������*��[�8]�Ă���$���[m'��4�:i��zP�$E�o�/�2&�������Х�'��:E��,�������l��H���g����=�*������3ܹ`J�`�5'���cD�rN�k`��[L�p��& �S�kV�g��� ]��^Xˠ�;�#��G����4;<��ߗ. ���\ 4W�	����2K�n��vd�L.��x�����e1lC�~	vjЦe'A>s�����%��X������	�+�`������S�8q�Ý~�tgc�܎묎�������[��?����OMu`���3�tߑ��v��۷M����}*�3��Z����K��n��9��d1��>6a����\���YZb�Y�閙�%�2��td*���%��p鈈Q/�����R�_j�HQ��%����k�`�Xo'�VͶ�Gn�;:�+kD�<=�̬�`Lj*���&➞~���lUW� ����4��������*�2����m�������vH��"
��UI!e�N�<"ȇوHq�^��UduW+}/	yo�C.A ��ل(AS�
���+���h���J���}�vCF�!ԓ�H�a�ޤ�;����HRS�уC7���rMC��a@F�,��@urzH��Z/�Ns�gK\ۇ˵�.v����/�4 n�pr&&��DP<�<�
�e���5FO���3UТW��U�~�m��� m`*������z�eˣ�g�>�GF�1	w����o���smJ�M��"�?o�u&T��2&�OؘT~_�=�>s�Lo��K)�<��{ӱk�baB ��TC{���o�B@}�ıi���@�FEa��Q V��ؓ��f`�G'&�LMQ�HOO���`���.�é����F͹�F���F)ju_6��4,P�<!A�e�2���m�Ȼq����4e�����%	MM �� �&�Qr�G:�ذژD�K��@G�ϝ�R�u�+@�#�i��b���Kf�f��M��[����=���q.Ȭ��z�y���9tU�d\ò��pi�xAj��-@�'ڟ'f�	������g#m>���J(�P�:��� '�p�bJ��$�9��v���I�(�����ųv�w�^w�77��1�(��Ǉ�������ՋY#r�J^� �����B*cTlB���
����7n����_�?�;oOM�
|8�ո�������BWM'2�bآ�l�C���+Ε���|�����H ؎������X;ݷx�.L���S.@-V{"L��!���+�ao愯i̹(ҋ����F���!T��z���<�l\U��?�� &	����7s�	�'[[[+�(�N���Kآ(9ݣ5n�|�����ݍ�F�o4nXё�̩�JJ�6�pL�I)����-﹠o���ѿ�ҋР�]w���]�oxx���΅b��w�Q��\`��5^�lu;�m�]��nr�������|g#u5���J�|��*7�\^�4	������ Ȳ��_�)��lO$�=�>��3�q$����������9��ZT�Z������^h�?�pV ��uϝc9f�铀IA�#�� �<J"_��"V�L{Է�o��6"t�A'z�#�}}j�Y4�&���,����Ö�Z�rLB�t�;��r�m��� ��4d�����>i ^d�{�}���H��!]E�Y���]�499���x���g�2�����H� t
y�f ������:��Z��3%"
�L�����>i�>�T����������5������I�����������T�Rl�i� �N���W�0 :�jjL [z�&! �Wt<�ӊ��M8�"m$����g}�@�d��N�?�:�	�2��p�~3�=K!�S4?����giee����wfQ޼u�Vi���l�3�Q^'�X�r��PN���F�ÁE՜�z��@h����v\ta�:��RaȐ�V��Ac���*�'��q�l�d���l����2�*�����}���J����(���dA�镑L�F��-u��	OX����,���ud%#�x
��s+b-'�tr7S)�O%V@i��,�3a�;�ĺ�S�����rCRGa�klW���$�5~|wY��o���}}��y8wI���P��e���;��o�,�7K�Z:n��D�UZ�Q�ܾ�|*7��1k ���@z�6 �'I���a�3��ˁ�p�0���56���|��	�G��f|�Ώ�3�;���s��}1*�sZ�䦘����rJ����F%��960|Ռ!�.��� \J�wv	��Gq�=B��ڕ��$i%+��#�����N�dR$
���JJ$��g]�?z����)o�����u�ou(&�u�����t��^(M�:���gֶ#��
dW��Cǃ�b��z&�������l���&i�����dɎ2��MQ��//XT�p�7�2�Ka�Q��4_���hblPmCCC����9e���t7��G ������A���;OЋW���X#ڎi�ǧ�J,��_?�V�<�D|�'�����v�x������/��� ��9����B�Gd��O�C��^���İÓ�k./��M<�8��w��yPp��`.��A;]�������dnY�fk�Z���-�tŭ�߻zX���j0;5;;�ے���vʺ�^��Zߘ�Y�e��b�b[���6���;�u�j||���3pq2h���<7%�Z,����籝����~��R�p��(txyŔ��C�j$j(����Q�t���Na�?�|NM���5_��U*:X��@�c�#7����{	�H5��T��������:i�M�����%{<ʒ\RU�a{�0jj)�,�*�^`�^�b�S�	������W�>�P������n���o�?�;5����G��l_�m�[���2��iii9Jf��])�ÈH{�S|ŵL"^�vtKZ����ﾱ�,?z#��揞�V xŗT�Sm1��r�+E���B��I�E�/�[�����.%���QLw����V��g�{�-�>�k ����=���;��^�cit3Ӽv=:j7�[���q��MVK��Q�I����*ݶU�w ��H�G��4�^K�Y �0�]��8J�z�kɪ)��6j�N�Rl�6�5��y曫Uf׿v�L���x6:4��Q��~������P}����Co��<�6~Jg���ĒF���/�?v����|U(K�����2"bʑ׻���cJ<�0!���fl|�+�I?��\rc��?*Fb��q�i8�iY:������q4ug��c �ɛ��g��PSQ���ճ�j������.1*.:J3���H��.�����%S�[�O��p��i�f�U���l\�������� ��p/p��6tHי�+��!F��9hu����x@G�T��ళw�5�� P(]��0�����6_x��XʞN�\V�:aX��|il��3�<}�ҨOyO�ak(K�`6:l�GZR�G3��(`���'q~�/ϰ,X�����n��Z�m��-�F�Cf'��i	��Q���g�����Z��PYM:������o�
a!���Xt%Ҍ�Y�R|
� � \�����D�_� �8�j�N��jt�迟M(!��S���cn�x��T��Y�V[3�[bƗ��R���^&~~����.���n�.��&���Y��ZM�e�q[�&gb�p_�z���{:��l�K�I�g�x_K�?w���4CÈ9LW�غx]��B-t��ז4�)��g��  T�II�@1sX�?�To���Կ�2���cOլ��$��U�&��e=v�5�K>;7H���~*�j��p᪴,n�o� ���w}:��YD(����J��Ƌu��l�*=�lښ�1q��&"��@B�͋�J�2{A KC w���U9�,9�X�$�����,���!���Ð�ȵ;�]��`O#�$�	\��oJ�	Uy����N��G��.�f�P6�GFy%4=>��_ez������E�m��K�KV�d�MnV������E���Ӎ��
��3�]w�:�g��d�Fv���7�d�+A��OfC�DD�z����ĸ� �`�xj�B��v�����H �O�BAv�zd1J�[�Ĉ�0�]�l�~���3F�0�H1��Ԯ���W{v��d�T�
�V�$#�M,,��d��(����lwƐ�*���Z#��������y�4�rؗg�ۣ~u:�۳�y�m]��2�`�z_��Ȃ��r�ni�����7J�Z�t���}����q���#~�z�:V�ʦ+�����3����
j@�c�t�r�o߾537��� R��'Q�Q��?��dLT
�opJV)rY��t����=�K�;ep4_¢C	rz�\���}e����1=u����V�����x͍�<�0j�:HH�D^�BaHj*�����A�r���7:���߶�$7�g��������=�=Ze�:Sy�j���h�s�(9hΣL�gJ��ͣ�K@��K�i���+���IBUm-0� I�<�Uʟ/�~Y�f���c0+�m}�ݵ��h���r��� �bQ���P�`h����&�72�_�6V�~��J�Z.#L������b!	Ck��?��7���T�Cub��ag���<>����Β�_�ڋ�|j;Q%��Q��lN/q��4S�^��������^ ���Z�^�|�H���䐇����	��@���8�����O�@��\1��_�֏7�q�p{�PH7�'����͍�Y�n�l��LF�����+���3�G6���c���#/�(0[���t���nZՊ.�՞@�Ej�Ɔ9	�5=@� p][+[cY>��B3�]����$!Ќ�h10m�1�T�c�OY�@A}�-1������^{+���|�j	���N��w����Qm��{�M��<��c�w�G�����������yCG��J+1%Xv�L�N�6p�����H�����>j��l��I�2P�_l!�G�zz�9u\��������)�r��`K@֪�+T_�$������#H=H��%C666�����*�ХeP�D	�xW��V�f��� }���ng�Y�Dic�8����� $M�x� ������ɂ�{�?�{�M����t�&'U�c:����JS�q�^�O�,x�#��
���h�������C���%�WX�6���{���s�Y�Θ쌊��:i.�ä������NJ$�HtX����q�*��>�NI�����6VH&1d���PRr�CrT�&��U�?5e��D�~#�|lm_�i݊�Z��x�A4�RU6�L��PLe�=M2Е�6]߀:W%e_5���ȼH�L����V�`+�:h�@�ϙ�vZ8�kk�Gal#��D�������.�?�?���� ��gӟ�����
�t�9��_�%1������9kʐ��ߞ��Bm��B����0P@H2�|�,��i��[�?o/�H���P����:��Th_�E*��H��:Gw��������l�
�fl/�c�����W>��~]�v�ӳ��>ߌ�
{���[q�~l�I�՛p�Շ�k�Bov�JP���4� Bh�;MO����������c�($����{D��������oo>���:�����#�1a��r�����M��G���8��`΁�U~|́�lp��)�q?C�cbf�jm-�r�IR5�����u�ad�1%xU���;���>< ���װ�)x�viG�5�P��ȗ��c�S�q����\�t_�_\���9v�9���$��	�7:��?�,�
ݖɍ;��UJF�Nu�](��-��'7{f�ֈ*�uI���yŤ`�c�/]@d�ԭ��[�h(
�ޖ`��`;�Mz�������xL�>z�ߎЭ0Hh>4��~7�qZ
	F������dx����Bm�ea�j��f�#��)�sU�?諔$u�H���py�b��
�ߧ� H���4R�a7�13$�(s���φ<g�;���Ҝi��@��F�·�'G2�K�Ee�aL�Vԫ��q�� 4���e$��ϴz�s?ap��!�&�ρ{�o%*ɗ�ڭ��qli�? 4�}�*�������[#in�9�D��)���n��li�{{0Zځ��s�֋_z��&�	ӟ�Hݲ�*��F��U���0}'�%%W[�y|��gKf�9G�Ht6P��`��{g�z���&75�8�.�H%e5hn�r�f���f�3i(���E�T�BW��#l����?4^�5��l���B��p��n1H<<����p 4���v�"w#0���4�7{>�1{�j���cs'��I�~��*�F�,m�А�Cԙ��u�Xp�C��
���jʓ����T��6xs�X� g�� О�4����X;oP����u~s���`ݲ����^�Y�c��@�y!���GP^�\rXF��B�+C0Ȝ[�)j�|�q/�ە'�%A o���I�g��Y��VU˴�`�%��%.��0ժl2h��P�R����ro�Qo&n�_+�}������U��G~�,����kzv��ȡL�?Ǡ���7�T�v�N�/�����&��j��p�Y�k/�7{�;�R�T�Y�rA��r�pp�Io:Ͼ2:�w���hm���A�BZͻ��a�Y���^_Ћ<-i��]���s{(س`Jn��P�B��~d�[i�Z��P���˞ж���q1���g�c��*gXQ��X�gϤ�2b� ���8�<B^Zp�iQ���4	N�|�5b�2Ijel�W��P҄����3a�hfP�NL�;��{�n"��f�ΤB-PE��V�ދ
��y�X-Y�l���ڎz�]N�7<���v�n�ta�ڃ�5���M+����&\i^,S� ч��`��C�Op����V�b|��7nXuL_���d���;���������_
�}`#������<OH��0�$�u|��$�Ўc��� <`��h��,�is�5��q�#����?��Gm䊊��F���W:Q�^�:[�`B�J�Vw�f�I�ƛJ̋�<W�ͤ�6e�{����{cƸQ��2��|�G��]����h��síp�DsD���ؾ�nw�՞����NZbؖHZ�v�W7&ڙ;wB˴-Tv�8�m�u���-VL&o�g=�":��+Z�
Y��$Q���cF���`=,�$��:_���(;C��%�6Y��B��%-�k�=z�}���~�%̹F�/6� �Z�d�ɬ\��?)O�����A&>u翃�����~D��>��Aƺu~�����ľ�6��e~���v�qJ�r�L�
҂Q؍�G3��`���ц���iK�|K�����w�����_�-��r�v=4��~Ŕg�1C�\j*�|=ެ���~�aB@�q�:�w�!�p��u�����Z1I�0��|q8T*�y!T�>n"��l���Uѷo.�c=F(�s�-�L�[�x����)L5e*��l"A��j���t�QE��ԑ��,�LQ�Ӆ����풆��w�6pn�_���!#"�.y��i�i���Fe/��,L��)�����Zef�a��M��?��$��.�?�p(p8�ej�=�V�t+��+�f�+ �����"�u�`�yM~�/[{��٢�]�^#��6�{�w����c��0JJ	�������qn��.���@}p�L�AV��O�g��4*�Ǿ*�� )9�G[?S���
c��ޯ1�ӨW&{��Z)�D(gH(1r|�(�^�<�����v*��4��j��i�F���\(����t�5��վj���$#�ԋs���@��&��������ٳ$�`N�%�`.Q
�d�VT������/�*�:��-�vۙ��K�f�X�/Gт���d����	 ��glI���uܯ��t���$�����X���r��,����L�4��u3g�kx���Y���57�{%O���@ӵ�W/&�(~���xv{���5<��PH�ۣ���GWA��C�8Ge�k�\C�̂&��v.��L����r�t�*�9<��3T��L��>{)"r	��$((�V9���~�z�P6�|D��菣��/P�12�Hb��T��s;3
�)�Wy]�G*��ٲz�&V��){^��z��g��t��sI��ή��I��V��-29��HN�6Ûq�(,�A���M��)JJր�Z#�H�9ߜ�}�n�IM��y�wc���[���/mWݯ����I����޴���y�vQqN_(i��Z��Y��]�����ۚ�G�D�\f L?Wv&��ɷ!��浉CEƵlW����/��B�:a\��}��D���|S7��0oO�����������B��7���h����V@�xp�;;�Vnۭ3�,--�	�$��:�ٞ�(�ѣ���~q�@�����~��(7�Ǧ?�T��� L�͎%����&;J�F!+�2%��e���LCs��gf�(�a��t�v�^Vgh�����9�MO�:����Pi£��q�m扖�ǳ�ǡ�����S_7�)��l��&r���"z���͆1��de��'5�2������.k�7~�@~7�t����j+5w�x��ߢ��O�lj��!��:eyڧ�7vN&9�ޛ���R����(`q(����D�M��aTk<uT�@�H��U��N�g'[F{@ª.Y���?��QO�Ƭn��gu��3a��r
Ғz�UVB�@��jo�$�l�����#:q,ܡ��+1IM�T��w��sQ�WY�����"䉖��gϤ���ذ�D@q�)�R��)>x�oK��"7$�tR�g㌽�*9�T�̥�����3�����=Ѣ���%K�__J�Go[ۛ���ѻ����N����;濩��sx��U�q�u����o d�d��֦�گ�M�G}eZiBJ�`v�W�*L�|8��\��⨵�������"==]�|���y������"��V�a��_���<��>~{�z%���]�:��%�����}�R�㝂���G�5�������U˴�v��>}J��s~��q����*����[N8����������G������5�ט�����*��š�����_E6��*S֝��8u~�G���#�3�P�y��p5��Ap�8��?Y���
��������z~�2#�"yE�{S}��2�{K�ǲ�������>U�����C�t�D����-a����Ɍ�-�/_>�=L��X-#�ksg���|T�k;L#�ʶ��`����E+2��tt�DO�����(�o
��a}_~�[M�	]��a~" #(��9�s!lޓN��ܝȲ%η-��a撓g2�@���{A4	JP0��r�d�YTՍ�/�����Wd,�o�v��Vzmc#�
�|�츛]П��:����WÏq�7UTx�K�S��?����S��$�I
��@A��h �\Π�!�����?���t�!�A70j���a�w�� ���=�<5�=ts�%Z�ps�wy����F���Z�N�
�^=?�Ӟ��y��m�����Q�iHA�r�<o�q,���7KsZ7&D`5�#]0չ��X;�_X��>��!�TzЋO#O{���d�{�C<w7�1�{*aK;����
�V2p-GY�s~ε��|�f�5Ϙe���=~���&P�ǜ�?�We6�!,W?/C�T�b]�C�h�%*B����-�O}7(#N�i�։�;=�R�ť��hAƀ�J�8����)���4�J�e;�R>�q��?6��)���ӥU0?���,%���O�e)C�.�fE� 4AD���5%�`0�`�=H��P�4F�jҏW���#<??�g��k��1���n"@3O�\3���TPv�hh�7G�2�.��Y�E�`"W�Ö#�'�װ�I�<� ���#?L��5Y�?r��T���u�җ{{�FPi0O�C4fD���ׯ�֟���2/pE�Zu�	-*'��?�
2�VJ߶3��WDA0�U�K5:����c��\���/>��=�a���P�p�)�o?��Xr8>���"Ab��ƾ�_��k��KɃ����N}��o�lm�o=s�`�,���-����L�Z�`��_���Iy��^z÷|9=f9}���8ս�!���a�Z�E&o�7��T�d�W����I������!+8���u
2��?����< VW�g�)��T	��v�פzm��!@U����o��-/@�+��4by��?%<����r��,��N4��jn������P�����~�oi��OA��{����k�k���g$�6�ms���R�#-�I�UZ��۞��=�Lh�B���m��yO=--�3�9�ޡ�Z�c��v��F�=�Y����K	����KBT�y�Ĭi.	D���0ϖqAǭ�g�2~':R�?���T7-�I��D�g	�	�~����m+�W�"�mmvgA���q�6$�Dr��ZA�lj?fE�<�_.	^���u<������
����z�e�Z@�+�mD��#��!u4��`�⒄L��뷁7���7<�,V&����쾇�[N>����l�~�+�urt���U�{�$t��:�ʒ�%�����ր����Jn��`ϰ�e6��w�~�.��pcm�a(���&�t^�_X�0Q��J2�R,f���+M��a��<b0��6wnp�z!ꈣ$#8�]�S��"���8��R���V��!�\�e;??jѻ㡷��=B��I��g�)L�����lYu�ė�Q����C�/!��ȡ��UHŒ�S�WJe�,����:2|Y�-, ����`����^��̞���c<
,�?
�D���g�^�^���w>��T��Oq�9�A���GK&5�i1����-�)��1���� ?w��� ��O�Yjh�0��#Tbej'�ݡ�'��;�|}�uR�l0����dxӵv,Xeraa9��L_�-V�;��m���jIɛ&w;D�/|��q�0�}����P ���[	�7�"W�F�k�-�7�FyW�ΎA.�Bl��ޚ-9P>����H(<�&spӵ��'�bϖ8s���#O�Ќ��Nq�[��O�hW�V"��]�p�p��N:NBd�5�e8���\t���gS�;ю�i�������Be�\��^����=�
�F?�!�9�ۦ�IھO��x!=����d�����M���k.���/q(l(u�hɊ��:'#a��㫎IOt�M��^|lllX��Y�5����Q:x�I?7�d�&����x�/���ux��U��u���\��҇#���qq8�Ӗ��e���G�k��˥��8'*zR�뇒c��}�/��y{��������&Ϲ;�
��y��.�\"�E��7��Kf�й4����2&+0C/�2~���єPB �H�H3����(g��U�![�c�[��M�d��(Zn��s�®�`��q�.�z�N"��&�v��/#
t�rU+�^K]F�o@b���M$���	Y㬀q�\^�N+���\��S+��_7l��`wWg�)�9�+�\f�I?͢�G�=�t�v�dB$���������\777�6s��>-
" �T�5r��}��m���U�������_O�w�5j�英��*�{��i�q�#t��F����8����Mb�I�Yȧz}��K��ѸNO�@-���j�̓M{+z�҅y�a%��Rd�ɤS"O5��t0Q{>(�d?wy����V�Mi��2�C�Ɋ�������v<��J�w�5,E������`��Sw�IF8<�z����`�(0͇}Χ�sf�ϝ�5V��"F��e���F���J�Σ�UJ�@�� �'�$,���[�����Vx��w�=�9	�[�c���CT~/ũ�1���5�3�0%�P���:J(�w{��&j�"��v�����#�L$0R���u���Ojld.��^�Ε���O��&��TU��z�����'�:ϝ����d�o�|�G%��D bV��*������1SOϴ~N��n�p�������-�,[�Jw�6���a��?֯�ă���ɠHp���+2S�XV<$y������FRD���	s��!�HS�"����Ic��<[��ju_Ҽ�b,�m��l��$�W�gk-��S����p����VT�΅ﳧ��ۣM͓��	׫��<I~�Ӎ�z�������Ht��4;7�Tx�S�Œ��3@��.��i����@a``��������-"Ǐ��$�	XS��S�B�߿,֙�TD����,�xTTT���,߳?���������'@ŧ�|�
g�)ڊ"fn�e>�+U�@����Zt���i�	���
��2�>�Z��,�[c5��~����(/����[�6�kƑ�(��2 �����P�5�{���4�����.�XZp��$�Bb!��&E��y��A�1ɗ����1�s>���y+r=�M����O�c�(�F\�P����5vi)���?W���]:5#�_�������d{��@q�#y��J�N��gg��g�EN[l:M�MF�l��ޠ���g/�l���=3gyJ�П2M��`����1X3��6���d�g~�'�,Z��`D"�O��-��J
�5�3�O-�Y�!~�0%��S*�[��o9��O�9��Z����#OO<u|�S�ɨ^L���P���	d��e��Y'1��������XV���IC�m�\�m$�O���SK�!���=!h����i��;'Ȭ��,�=���A` ]����ܡ�s�+d/fޟ�V8��3T��(Z#A��F2ɕ�}��LP��)���jϾ3y��EA4�ÿ!�I|~��}�rX��V4�=��=1Z�>خ�?|��f�f�.��m������Ӏ@�N�.�M7��xAZH56qJ�e��a��MNid�lw~	u�����`�����T5���л��k�И�������_�6< ��p�)�����N{?\o�p�C����� (�o�ě�)I���Qr?V��d1�)kO�qC�>D򥢽]�:`�^�*Xt\'7�2{4r{I�����_[÷�o�#)�#�Rc��!��sl]�Ti�1��_�҄���P�����)����n�sc�|SU����������ܗ�4�	�t�=��"1���m��)�	���l��Q���F?��Fkw���O��O.��pqN�G[O�gm͔���KҪ���Hvσ����Z�Oϩͧ�p~U��_���{��J�Jq2d��~�6��p��@�*���F7�iQ�`ۭA��8[�� r�#Mg4H��@��XѶ>&��>��(�S�ߣ�!(�ku!|��.��k���?�jQ�(�sE��\�]�ׁH��������c("Z���G�G�:q����C��v�����0'p�3kR�LmQy)�u�&}RU�h��)��;X��;2��� �SQa�p�I��l��x���Ã��k��QMM��k�_嶭���r�J>9@�bs�#����n�8��3�xZ���_�>=�����C��Y@���o�\�Ve�X���w65E���}�g@��� K���^�r�\�ZJC~z�O�� -DϞ5@H��K��D�l��\�zX1���&��CG����ƠT��y�޽����{�{���˘������''���>��f������jW�^E�^��˨V�q���,�l�ZM�y��XZZ���
*�
j���c���ݣ(�ds�ztt4�����7��f7X�B�=��h��]k�eo�M��,K��Ǐ���L�|]��0133�ջZ��̙3سgfff��".��ٳ�/i�F%ۇ9SƵk�2���O��(�3g�qN�N�s�ضoߎ��%,,,�ҥK�w�����T*���֭[�s�N�B�lf����)h�q���4C���ܹ�z��z����E\�x̌������:-�8���(�Y}�"�=�!2ײt���2�og(�� ���Y?~�����_<|��J}��F�W�+�2����f�����>f���oI��i!��9�{���"�ipY���������	���s�d��!8���&�A�)~�3/��h��-�f�N,�P�a^3�܀��̏�N]���o�4�}.K�Y�׳��Տ�U��\��n�u>͠2��777�����>������ݻ�W�7C%$I�Y���H!��I��_��������D�·�p}��#_k�~}&��F^����}������m�=�&02�M/x�e��~ԹW���g~�}�/���o��C��D����+��P*M���{��O���i��1��Z�}���ر����������7�[�g�f�9��zx����^�7�ٸ�|w-�� v�����a����Z�M� 6���޿�9ڊ���1���7l��봙~l��4y_�A��ߑ$�����v��ѭr���)���
?��t���?��?�g�<p������o����A��`@�����GSSS۝��)��3�^��0��g�~1�X,n�i}��$x���c�Q������ǯ������2�ES�ibb��U9�@�ݻ�������(S�����Mp�����H�ػD� &"-"Ph�) �Ҹ J�G2�̬ P��-DQ��0H.����:"��RA=�S։�	@���,B*�[f ���v8�Ի��>�vu�F��o���G��ז1�ވ=  |��NXk�*��
�P�I�:�����6#	H� l"�Oi#%Z燄J 3�Ŧ�[!!2V�b�P��Dƈ� B��rf�B�H$![�u��"Rld)�I����zL*�xJ��k���� ���$Pd{�'�Y$��rb��Ɛ1�����K��r�M��dD�0��T��0�a���lL1SpZ/"!bÜ:�ot:SF�<3�|~�K2ݸ[&+6̅_�7:_��^@m")��(�b���2q��`��Doa@K7�d�D4��N&(0C��@��C)��� h�:M�� TJYf�"�Ř6�z$��Dj���B)Cƒe"%�F: e���5�%	��DZ�\E=P�̖�%
z�w�Ek��~�7zI��0zcPD��zgV�:��ט���F�D�fٲm��S[}|���A׉�E��-=���D��d`ź<�@�!�Y1�LzM�"C"J������Y+L$���T�e�$}�D �DqZj#
 �E� J"���A
�b�2E�$ʊ�$�6&k��E�Jk#�Z�Z��*�tq��Y�~E�;���- DQ�,IL�Y$
�c-u���֚����2i����DDʥ�}"
ED($bf H�a��	��Jqgnn��(������9kmh�i��(��ur B�#;:��8���~%t���8ON�(ȋ�    IEND�B`�PK   �cU����:  ;  /   images/71057ff1-f3c2-49c6-8a17-bf9e68e09ed9.png�Ww%��.����y뭽�m{�momۺ�����m�����wΙL2�3əL2y�P�#B@@��H���'���'x���A+&������z�������(D],һ�sWJrjd�!���v�:a���2�	�Mh�~L&�X��tF�,f1�*8�⓪��UR�	������I{��
F��E��A��s�w���D���H�-�>9=}~{���O�<�V���f�}���./����?>|���_���ƶa$<��WvN����~c(���p%{�&�$�f�g�d�������K��˫*+jkj�kk�s
k���%�=�cc�;[[wwwO�O���[[�����}CS��k�kmm�N��A����Ʀ������ޮ�����CÃC333���Y��q�	����`�?���2*;�z���@aс�A1���IIii��ᇻۭMMC��[�K'��g'��S���==E���Wg�w�O75e��Ԩ�����x{��8fe�KINn��-��sptJOI)��365��kic7>2lbfVRX���k`h`ni��������P_�1����������)((JJIs�񋋋��������*��/~d�)�'�]UT����$�Fp��r��@��C;�M! ��e�E�<�/�^V��{t��ꘫ|�{ל;�ҭdA�<�ۋ��X"��
8��a�n�T������WlO��[OX���6>|5KO�^S����^G�}�4�P�Mn����5���:B��e��6��3�����[�� ����D�*�a+�Q4�܀UU�͏�8�����<b���_:��nΥ����f��K|��ɤ�j���'v��gm��%!�)��:zz�	��Ksёeg�'Gj
����힍��|B�%�j��A�W���n���k���{7z� 6`6�XJ���\�� ��͎��]����@Y�;��a��أ3�O�&}��L�Q����:Ut��ߒld
�"a磞��]��>5�_�EVX��5I�k[�8��8��L����R�����W�h�kik���s�U���<�#[`-h�c�Uw��fh�tX��!>$~������'��|�n6Xڄ$�泫��H��Oq��0��ʓ�V���
�ﲘ^u���������^�s�0���`
ۮH(S/�oW�X>:��k�w�Px̧���٢�d��:�^�^��X�8�Ej�J�O�ء�펊�VO���ޚ��<z~w�K+E���V�D4��4�$����u�C�g�։�.��^�*
;v6�|P�c�oM����|��>�#����W_0��
���y���xzy���Pa������F�)�����p�f���ꮷ���|l.\��
����H�Z]���/�����W���cɐ3oX1e�n�1�S��l�Z�S4��6���Q?EU=>��)��	� 7"���{QM���7W�Ĵ�y��a�~b�_&��9��i�Vf2'۫�t_Ǥ��V���Op�2�+�g�K�i�j��Ó�U����v��ڤ����Nnf��]^��`�&���Ǧh_������zMͥ�7��Y��͉?(�v�z�^w��U��,4#�j����J%�0��O���z�!9��)��'���I�=<RT�4Ź��~���&���a����=�ޟ����ϻ�짜p��p�^�9�6M|�J������W��51�-�.�ױ�>�e�O���7L��e���߭������ϼ���o�G�-�?�Ǽ�4�R����r%g��/�71���{�.ef<mZ�(�ݞ6�چ��8�'&W|�r��s�@�^�/�:[N��]�<�=/�W�f>���F����ĝn{
������_46�*���������ᦦ� ����k�=L�J%]ם	���V�Vo��Hv��n����P�^��U�s.�8���#
�� bjV-@#�c��!��M8���z_#���u;�n4�45m\,$��)ŧ��1t��C�vksn+�r����'	�1ކ͓]\ ����[�.����I7K2�_r$B�`(��7H#��@:��?�6k�
����JZpU� ������42^�sn{�V
�%�KK�3K���Pn���M+Iu� R�I�6��v���Ggc���cmO���i��2#�	�EC2N���KEI�b�٣�7R�y������>��#��gl#R�1-\V�&�L� �m
/�����i>�5�]��Z�}j��������4kd�M׵<˝�R���;�����IGWT�癒����'���v�m��k�}��T�F/�a�?�m��g�a��������#+̺�$�������Y�}O����~*�=����7�q\��K�������<>=w���������,!���t.�qշ��ԥ�
$rz�2��e�Ҍv: ���T�%���=u�E�E�</RＯa��$f����.sE�C���{����K��فA�s��ǉ�X��q�L���t�Z��DY��dP���"���vJ��pnqD"��b~��%��&Jx-���}9�[6_)a�z8�)bJ�[���� ����?��7XK����:~c}��1G9q�"��g+�?g�s=Oq��\�w!�=�I�#g�
����zZ6�3��]<����W��~f�i/f��m}t�/��� ��<���W��t=b	q��`���M�G��9����fC��3��]�-\��$�Te���Sv	��u��:����ʝ_�)��X�\^zE���.7� �Z�o�{�b��w���TT
�V��[�CO �+@��~@䌥Q�}�\��ɽKF��tA��s0^�À�r�T�稝�g��f���η���]d-�#=ҷ��8c,:	Z5�i1Q摃yK�L��<S�eI�yKg�j����j�㪝)�$�Xkۛ�2(�TB�|�
X�b>뫷��2�ʱobm�;k��	�̔�ō�����
�s�iz�bc���+�NBܙ�tЅ��L�Us3�J߬�;e/Η�~��f�S�F���
�M%��4��$��h��G���?I��_�\LYC�����oD�C��F�K�BX����fn;`U����������M���|s-���)W�(˶�nA޻���?�ଢ଼�|���$-
N��aa�W�4�ku��"F�,x�qٲϲ8�h+�5�&ў�fPiO�5DC���w���7��Uxb��\�e7��%�O��?AO:6�a�>�e� Ioh��F1uq7`�D�1N"��t_j5���B�@@��m����!��\c5p��[�%�V]����}�l�<��a]��a[+�ag�I��m���Y�7+��ʷ٫L]���<�l��\��+��O��f#���ǡ���7�XӨ�z��������w��c�H.�acb#��%{�5h#�ݦ#
c�L�H}�)ș��j�B9���£D��ϩ�(������&$�¾�r�3������*��_B#��	��q1�\��!�H\��Y@����,��)���S��HPü��"��-E�!h5��a�c�^a�M]}O8@u���Uk��ͽ&��U&>.;z,#4�0:捓�ʢ����C�oκd�&�i#}!�Y$#��C�+"�]TfV:��F�`�F�i����zӅ��%b~��c���K���{e-��M�=i��8�p�7�ղ`��=���5���;��'�[�˘�N/r�I��x7ΰ\q.k���;t���T�	�k5*�`-�~������`%1UU?=1��Y)���Q���J�qr� XX`��8�c�{�د�����O���<d���dx��Ls�.Q1_u�w������x-ހy&�/�\���AҮ�5]*��wI�˴?���`���X;Es�K�4iɦ=7��3����}&t�)��ꃰ�q������!kh��:eO,��*�i=�ݍ��j8↹��)��������!�R:�R�����-
��w��;l�Սx鬠,Cj]2�P�� _!�Б(�o.z��]p z�*��~l�$�2�N���cgqG�Q��(HI�M֭������s_)��$Bk���H1�2���o�
?���������M%پ!���(��E�A=�"�/ +2�`��r�c⤟�/Lm��&
��mco�R���x��5�چ���yz�5m�KWD�pj�,?Z!�a���$�V����ѓ��1�ո���L������ �\@�##��n�$*��q� �Y_˰���nQŇ;�P�.��N��^Z���;H�wx|����RYN�a�0��*���ޖ�Pt��%X��ug$*��ֻ�I��ރ��7MY�qx/,֋9��ٚ�-3%���1��!p�J���ji���֮��؍\i]�������qL�{�
�hy$b�i)>b�˞������I4`��E��e:؋�C��W�ِ3�g.�ϴG��c�|�7�FΘ�wu"���u��*�����-#�*kզ�x�y5h<��0b4�N�����4רI���N޸���!�}���/򿇾���_B}��
&+O)@��ܻ�Z��@C����3�1�����x珜���t�
m��5B��3ua��H�� rW��߰m�)�4_�K* ���h��F 5��̍赜����,>�+��_u��Õ���(e��K����e�Q4�2,�69��#ZA�Sm�T�º"�b#��F�&w,�4+�n��[�;��R����"7, ��!y����Ni�(����d�� [^�1�:V�`�
/�U���#A����ZD��Q��ɯH��fe<��q�w&s��Eͮ�$|�h��x&Ay��6o���BZ=��Wlؾ���q�� thG��P@f�/O������,��0�w\�/hf�=Y�����\�%=M�.�g	n���[U�;�UK�P$� !��=W��9��Q�=>��i�E���%�c�n��:��m
�0⦴�cU�h=g��^�+V� #WA������|*I}��M*�a�z󞬱�F��s,m|?x�b�σ���x��y.R7")�z��{㘖;5��`��`����10S>_�^:Au�g�������<�k���eliV��|�����h��rlo}w[O@�O��)��A�02ΰn����$�a#�>%�+�#Z^`/�	\� `����	%:�'te ��L��n�ަ�m��hAI�N�(�8�����2���~��t{�]�I�[�I�� - ��u��JY�HLB/�`%���c�G�Ҙ��i��_#S��`>�Bӹj�ʫ}KQL>����g*�G���b��$�`�]Q�,X;�;B-�)+�Q}���`�OXB��|4�T��OE�����UOA[��1k��S���.<)�,-��dF�֔�ĩԠ� `Y�b^�����@��u�������x�o�ۏZ��(�*RwD�t�����aBP	�?Qx(ưx���R�pɒ"���SQ\PS��P3�8��a�\h��sQ�5|J�.�	'{D�F����q�ƈ+���֎F�b\�P�*c�����A�0Z�`���ʡ�u��"��/�p�#��[�Q	=W��E[�����/������$�+�h�X�D�]���q��$ `hPE�/vY.Ҧ����\�����i��t����|T�
k��.cpBA��𼎘rM�;�{��/�ŬI��T�Ȃ;�B� W���ڨ[�e���?�(�N�E���E�Tf!�����2�{��$��f��p�`# d�7<�,��S`4�-�q����o��Kg���M ���2'���������*���U'!XAGVT�vBjdw�"=��ϝ5�i9�p�F8M���2r`tp��Q[Ou�����opv�i���{��� ��<E<����()v�:@��|pϿ߶:��qǁ2&��m�b�X�<�6�h��P����7�&2��b&S�Y+~�	rۍ0�P^�#p����=|�\�T#�0�HQ+]��ң�0q����۝K��4e#J�ե����=�t��'@�&�(
��>�\+�y��8�vn��y�e�����_d�ڏ�
h5���o;�jk�@��g#�wo��/tm�C9j:K�Bt�ɂ*F������j[k�L�7ɺ�~[�>��}J��7��`;���xsb��0T�p�T��뤣R6�=��)�����S���l��AH�6Om ��
{]o\�ag
��u[�?�d��+x#^�	�P�5�<��q�2h��?�'�3��L�ԋĨ�%p��u��1sV�C{�\-�����*	1�	+����ۘ�JȽa�x���}��F�"��Aaa����q�`�!�B��\����ZX.0x�EVV������#��b{B3q�$#u,����w�^��Cb��v#~y���y�Lq�B�5�J�uriLH�=�彼V|Oqb��7i?$O����z�Sꡲ�AK���6
��҄|����F�:ݼ�'Y{�n�gH�=3
���H��Q��g�]�m�t*4�̄z��"#�ͽh�U�W��G$㾶C�t)�zK�������z�Q�D͘�:E�����b��e�ŋ���2D�6Rޜ�J�H>�!�}�������f�o����&���↖�rq�}W3�ק���wz���A���X|B���L|��:�91�����n��(
[�d �]�@�e��~:Y�xf}P�#�7)�h�X�o�xn�'`��>bP��$$�H�l�H�B���S�����S�a��l.7��~��?9f�� f?4�P�[��(�;<��#���(�*�$V�cƶM���L?�=�8��R�#�'H[Ab�ŭ��͏��Z����=T�/�����/ (��ZM�/<�_L����}" @���5>���O<�ʸ�aQ/#���!˘�Ĭ��B��m\���p0M6-ǀ���in̠�e%w��0CV�y�Y��j��t��HK!	��<�/����.C�����N�od$pJ{&��lD�E�n��qa�F�ia�muE�Űw��Hv�ɱ����� �@������3�ᡕH�I%%vr���#ٽ7�����+�(���h6�h��5 �`?��9�OI����!��Y���k^�%��Z��n2U�ݤ�h���J�R;�qwD3p,��X��
5F�'}6+�/Hu͸�̠������E
�ǣ�������jŕCY��VA%�<m3!���%;�:Q�)d�����MO�2�b��o�l|>�H�Z<��C�q��˅a(*L���Rv�c��c������@K���Zʸ�) �/]�����`P�Z� ��$�}���FU/g���޲��E��B���7. ��hm!+��O�6	�?$vLh"A�%�?Q��'�#(�gqG�Z7Ha�:�ߌ���y�,K��=�e�߫u{��4ܤ���@n�'����N����˨����7�����N��D��,0��04��3ӳj|4T�������5i����$RZ�M\��$ws}�dyl�I����(<�J���J��{`�`��A'���$ɿ�(�~�Az�<{v��uQ+�[����&�*�+�{�l��8�������1޽حssU�Q6)��#@��������I�k^?d�4�&�\�)n�g*�N��E���8FYJ��Cu��$��"F.��<s=
�%NBN�G��Q�
�����OI�h��e��G����;<��U�&{�+R �8U1����UFx�QQ�#�,1�:�j�L	w��UPH;����ɐ!@d���5@�4m�2�W������ E�����_W�tE���ў���A���Н�@��}q�1<����a�[�1���Fȋ�����m�X��E%�Z�����@�q�_4�|�2�8%Q�������O��yP�n��;ڿ#���k��'w�A��@�cj�xu
L|�R�R��H���x1c�G��8<uf���@�)T�+P���,�m1|�L�"���[�m�k���}ê{=eG z�o�{�t ��� HJq��^��=Rle Ob	.)�QCtED�2�ԩ�ZJ�#W���N��v��j��O����*�[~�����u�̿%J6`��$�$[X�~ݷRmsK而�E�&ܑS\ei[���0�P�Mq?��<c��h=�B9r�U��UW�\OYl�Jj��8���PSd�U�L�ZkL�A��j}�c��+�0�`R>1���8��88Gyp$�מ��cW;@�h��o��-���������$�v�~�+�f�:�h��%SH{���^C�'>"z�/�����ʎy:��22(Fd+��qJ�⮉��1qأ������uYDJm�-}"���#�������X���o#f�&?E�m7/�L��5���v� �>�α�:ko"E� ��w~�mX&���}��ə} ���ܸ}�B�0f�,�Bг���x��!x�@���ܓ␟����/�"��z7�2S�F�D�5�T�A�w�X�1 �K�3����o#A���0�y$}c٢��29��흆NzU��ؽ�����,(�)���ha�b1k�&G�M��q�4{1fN<�@׫� �K2)����Q�GS+
0oE�n̞�J������a�c�D��ii�m������b;�C�琎��n|p�
���X���2����%��2�!�t�������T|�y)�d�6�;Ѽ�c"�h^	�^�q�.^�dv�f�3��A>����kEl��E�~^�����.��֒V�	�����7%��-�����E�h	��]ʨY��{��1�"�E�L�Er@������% �hܨ�����娢���;��(�'���ʆ{~52J86LŒ$V�W%��.�-8Q6tdk3G�H���|՘(�WM����k?l�xGr���oAF�hf�����v2���ca�$'k}U-c
a��>{�,2?)��b8
MT( �"���xۺ�z�~�8cq�߭H��[����?F�򟹦ӝ���6��d���n�����������|�7v��ϔ�-�D9iy�a��b�a*�u��XFL�@�������5:pIt��(gm�CG����ruQ�,��WbK��	�A�a�u���t�v��R �P�*�C���n�j3�YK&�� ����C��V���A������lRش�4�Q 1ׇ�@Ac�4*�~�0؀��٭����:��v��S��Õ���}���&Ⱥ��S�LOFJ�`ֈm8΢=yl'$�L�k��C�֜,&�=BsțKEU�l~�N � �&� ��a�w�{���=�Xm��ĸ<:��e�ܽ���r��$�ǽ��²��5(io�ȁ�����}qS$R>�8�͈���q�i�x���@r�h���b?xK�B��y��٠�(%���<y�(����Y���fÙ�"�fw��qӱ>�$Q��|�Y�Z<��ߨ���%���8uC\��s�36m;��HJ�gF�n1GX���Y�{6 -!�`����?�SM�ukHA��(�0#ޡT��VUE��F��HR����X�����b��jP�|����MU1ٚ}��ǆ�������]�`����6�(S��fb;�K��N3�,Pgq���y�F��&A�-}��0b����\HI����8 w̄!X�z��Of;r%���zK��o���E��F��8B��V��XZ��x�V�<u6'�OqIL�̖��#�"'�'��{�d�
�nB$Q	�.y{���#:5"fO�܉?��X	z�7��%���c%�N�C
���FM���P��.4�-f�R΅�=M�K��%�{���p�}����P�.n���3!l��L��T�E�d�`z��1�t�v7qqYd�$�ϕς'(y,E�rl�+z̀>sm~'I��O��4%'q鸣�������4�+��p(x!O#ה7�X�&3���� ɢ��Tb�L	˧􁻙j�s{�B)R�eUf�@t���O�8�u�����wD��q+��nB���ܩ5��V��׿v��qw� x�`n-�Pv�u	!PKb��!L�d��߅�$����<i%�'�>.��`v�fn�n�(C�����Hc��FS�~Tl}�x1��ǐ=c�]ɡؾ;�w,�ʯ����j8��	�U��X{���b#L�1�'>	p���4_��=<E�G��%J��o�s���EG��l�ȹh������r�p�ȍy���'A�v�X�P�T�gK]�o��
dc����찥�eޗr�����Y��#�KB��*z�|����ђ��\�ђb�����i�R��c��<���Wx<F(���%1�7;��o��ћ����{^^s�����D���Y����L7�<�(��xvl<�"Q~��}sY>p���U�@��C�'[~�B��'oc��Y�ϔwҘ�k] �l���1�懡���sqgH�h]ޓ�8Y�ۺ��b��"c�)��-]g�B7��礒v�
�F$d�� /-���7 �]x��S{�H�t�^H��0�������4&��Q#�t3ָ+ч�Iۼ��'�HT�`T02ڊ���>k�*y.E.
�����P���$���&���_fx"P��m|!�/,�q�G�k��W-�� �e��i���Vd�N.�0��ꦹ��˰^���X�ǔ����1���H��V�4C$f��gD�4�9i��i���<�[�C jz�"���!((>�j�oN��C��9���v��U�i���_%���6�>���^�$Zo�qv����oƎ,����zIP�ʥbc n�P	 W�F�c����>�zW�T6e.A�^/�Z��ա�0�Da�C�?c��ܰL2�5���rK�4�S۔�r0��wy�k��i����"_|}=��DA�6gN�ɿVA�����?�<1\+/*�����`, M'��B��8�C�2FI�i���Q��/j��p.:�}}M�熯���NyҊ+�|��Rݳ���Ƨ���[�V�D�)�na&K��f'���i�i�5�1�+��*���^E�^Ͽ���D`��~��4�@�h(ʯ$'j3��K�{�Q��+s�;���$<�6xm%Š���˵����@�i�o��xe�;����v�}*]�>ՑZvqq�8Q62JP�)����XU~ E5�m�u��5�T�&�ԕvѥ{�a�~Ǖ�l�P�K$��U��� �$�^�[��0�������:�r\���x�N���������ĥ�+r@�9��V����M���;{3��.���y�O�/+��2388Y�!����_�?%�<�y�~�(���u]=�n������%y9��h,�F*v?���D�燋��tѩ�������*���<�w��Yx��_����}-�\K,
���	�J&�ˬ(d����튧WN�;g%%����7��}-�tikki����5��B� �8�n��Vp;�qo�b��{d#y���dD!����:�ֿ��6D3ϖށ����v�ߏ�7���L�O�������;�$��4SRSFB���6���#�ڽ\f)��h�dWJ�ԖMdU}T�:�ǚЪo4���OV�8v��i�wF3c�Ɋ���^�j�?��i��ENo �1����������j�[�&cq�����#K������nc�[~�헒��֯hzh���~W���aiG���	peۅ8E{������煃���������Z��= #έ���{K2�'dkw�wA)���j�A�������˩Wx���J��Sd��VM�괧i��ܕ#-�.���B�	�s��><<��Y�@����hV��U��K��d��P��P��'ԭY����\'��>�)!b�t�(��sJxwwt�cm�;K����B��"�<�s��IT/]F,��.�XH`$�0�E���n��*Spxa�td����63�G��e��[h���"?M��
�z�5��l�ԛ.�#�N�b�;Z��[�7�D�o�v��ˎ���=�#eqzj[لJӻ�5һ�������4ԓ�[f:��%���yk��%�&�ӘWL\Љn.��#�s�>�*�*\ B���80�P�Y��#���c���A������{i�S�E�0��I&�����������>���݈���+��
��	�%�zu�m&�Lf`$<N��X{��d�Cʼ ����FU��Rs��\�����ߧ�A1����_�s`2g���~SZ��>~@��~�,4l�ᢈ�K���F�K���������W���07�r��W�O����~�5>��m��ܩ���E��p�x;�����i�����C��ǃ�6�P�����+�H��q������y��Z�h��V=uO�2Xx�:��(̥!�(&�Ք��v���N���r�,��Q3���|̻���s��ơ�Y����S%��)�	3�K���ي#HC��f{�#�A궧ƀ��2Z?V�ݴKunƥ��[���ڿ�an�_ �������Ƶ"@l.C�u�đ�NXී]2[+̓.G~:	�˫����J$M^�*�O0;�#Ô5�㞵�cȻǁ���d��w[%�[��v�27�}Lv�1����~�����$zyMϢ��N�����ڊ�����6j�߿;�͓��ݑK�	��I6�/7�s<����v�R�A���uu�99$/S˿��4`�S�;�۰����r�̃�緼��C��	b,kKe��|�2���>�Ż:*nEJ��	g��<A!ӳ��L3.q
vQ���󗆼_SR)�ܧƮ��y��	������ήq��_z�m�:��ܿ9�}q#l����#�d�c��Y���}Ir(�����+�|�`�1^w��M�j�t���7A��:�f�+[�q�˯#�� ä�)�J�7~��ܑ����ݠ���U?M�b}nc���Opc�y)�e+9�>�	��CE#Nb������l�3v���h=��)-�����f��ih��h]0z�}��V�h=Z�|E"aQ 5S|&Y�(�P�{���p��1d
���
��o�H9�:�]4/,psҔN&����R�n&�z�;|Y���\����	��>{	���e ��J�X��h���r���K���R}��+�P�����N镥��Cg"Ӿ$���iM#������c��{Z�`)��e���J��3M����5v����M����fy9z��^�#��
'�^�<��"བ��Ĭϩ}r���P1-ҭ�O$�_�n{Gյ+���q����c�twj��u�ܵ�r��:�Νy_-����i�J�;U���t��ڿ�&x�5܉B����ǵ�U�x}�O��� ��c�*�\�2=��d3�������\j��O$xqg��-����z]���&�ާ1��E�3��&Dr�?�8��V�wr�__���=�.�>:�7 �T�~���eih&@n'½H��m����Q6�U\�n������X��{-�R~7De�DM����Zm[�w�0���Q\Rs�s�T��fb��[�^Tu������KXe2��Օ��t�����v�'mT7��&��lm��[�	��٦5�9����\�,���E���M퀔<�_��[���N���4J��%OR�Q���-�h�١��#��O�J(�	��{�WϿ�&}�&;�w�P)�+��c�CB�
( ��K|=��~���#3�ͽ�����c�B��$�;��2
Zl�����L�?� B�U��k��X����m��(�*$��(\�<�S����q��<r�l�����B��t�J����Yj�4�EgF���ճO[�C��0�#��=��N�F��/8�u��S�I^OmW(�n]�+T@���ڽ�z^�F�0�"Z����ؚ�|/��.�Q�o���&;����6�n[ϋ(�������o8p��z�W��o��>���#W�tf�����m.*�ᴘRC��p9�Vl�rpH	O�E��s��ѶRoNZ5���X��]�Wt�#<����f�3b��+ʫ_Wq.įW�UJN[=ȩn�j���.=U���8�g?$�P����<�O4]pnJ#�h��r�u�nuؑ3�#�����d>)_=<6|n�e�V�=>�D�=��vq�/t�r�^��|G,��~J����yh*"�Ū�z;(]�����Ȫ1{�:2L_Z]�f���� �#t��+{��(?����onY_}�w�x%;e5��S6�?�6�.���9E�w�rp߯	v!�6�<_q���xƚ�B\�]�xR�������%}:�����t��J�q��*�ZQ&ؗ��O�v��}ܣH�4�����Xox6J�3���_:����AaʡCз�2�l4�s�����2�>��U����i^=����,o���`?N�u����f�$��3W[a�����]F 7bs�&v�˳��2X��������s�C�,�T����m��vQ�EfrpC({��[��~y�8���� �Q�%s@n���h)�hVC�H�g�v
f�{�o`��� ��i�,��!��^��
�f�߿<���R�l9�N������:�NY�·$��,�?�*�R�`��n�8���_���/(r%�nW�J��8QK�Ch~L�lW�{\��o����؊�`��F���"�[������,;v��S8�*C��#����Q�4��Y��H�-l �WH�JCH5W���$(�����Iv��.zl�4=|���$��� �_����F��u���I;B����s�^�W���s�9!�#	�j�a��PK   �cU��g� s� /   images/d4dd056e-e2cb-4614-accb-0aa130e74534.png "@ݿ�PNG

   IHDR  �  C   ��]   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���|[z�~Uus���^��uj�JD��d�a�͌��0�,A{��<˳l33�����`[�h	�n�:��{����s�9�[�Vխ����]��e	l�X�s�s�>����oq�S�t:���J%��n��q���8i����D�V���PG�:@���[���<x+�+�*�dݻ��2x���i�:�����K��t�n\q_�Y-I���=x<�������?=������ϾM]�\5����GםvQ>
�W��(�F���9���Z�C1X���N����/�[��ߦ��T�z�W O��L�*��Uޛ�_^F�3y�ыz�JF=�|��8J)7��G�/��?��7���>���z�x�e������e/a���2�.* �K�K*��?|����4��R8K��a-8ᦗQF��{LR����x��{�/������'Ͻ<��;��a}C曎w���#�U�]u�:��-����$��r�t�9�p��A^=<g�޳r��Rɡw��}����!S���-��z�?�{�����z���=�#��y_#)듙�t�N�)����BISp�&�V}3_+�ܿLTR��F(mW�1?�u��Rv�I�!�����}8��k�j��߽���Vr,W��o��R���͵xicK�޷{rd �b�f��w3_/
.�Դ�X�ʵx)r���K���\�T�M���NǨ���+�d�P鵁yy��?���zp-��C��{:}�3/��$'
<��|�FI�{�+�̃�U3�L��>q�;��}��������r/���(��>��B��4Ik^V��_ �5��i��J���Z�f����C3Q����Zy ��z>f%%�Rp;G��IV������'���gTa���"E��DW9x�g6��ȒJyV�@a�a�,�z�{}(m����y&��t:�^? b�'��͙��k�46����<���\Q/��o�۸�l��%�S�r-��F�s�'��3!6� �N��x�.32+k%�^��qE^�~<�|�{��ˏѽ_-���J;
_�|���<H�� ���ݦ=}�6!����X�,�d�e$�g�w��^�V`���<��fޥ�=L���VZ��� X/��RaH����\�o��<���;`I�#/�%��ц�[�W;�|<[�!k-�C�:P���5\��
J��c����@�l�����ڼ-��LlyTB�O�n� 0�O2��"#�
8���Yr��z .'=�Z'�h�׉����mf>��.2�v$���&.|��S9�[����j���H"7Lʑ4k �I��{�b���k��I��8�c�tVW-�ͳ�M��*)o|�t5:x'��:I�|��n�c=�8Y �����J>��	)�����4�o�s~�f�N��Ec�[!�%�4	*�fq��
�I����� �v�:
��6�8��f���-blXH��l���`�iG�"�ɻ�F�������.�>�~��}��	� ��=M�X �׭\�7'ʴ��_$�Y�w;�rMk����W���HOBKP���׷���zT{T�,�ʒy���c�1E�H�>�t�N��  �}��S>%a!��*��(�?�ϊ  ��)�y��	�ꑁ�@����*�4�DNEmP��Uv2�0�$B�"T[�\ԍ�!��"h�C�dfYW��@����-/)Ńt�VEX(�!�T,�S���I!"aZV��̓`���q��z֓*1B�C��	i��pt҆�JYEy���y�ͻd�H�i�0���ͪ�%�HRy'��+�k ��XV�ɋ-�GB�5i@���$~񘹶�ȏ�m_�!��B=���A��Ł�!��OҞ��`�4�?�����ڱ��*��,�@0/��0mg�X����@�Y�·OiU�o�=@~
2��g@i��͆��*+���Rz���Ղ�6<������"�.0�n�{l���W�Z��$�c` ���$m��/n�0����hAK-��K��{¢ĆG:�L�_��@���^�9�����7�" 3-8�r�J�2�T�\f^�fӖ�D���mf$x �2��'���0!�tI�d��	�h^Ӿ�I��1�|�b�Z����2��׀_�U��}v�h��v��Q�3�`�6&FF1ܠ��{`(�I�0�ć�B�䔲`�'����=�թSS�|)����OdB�(�( ���a6� � O�w�d�ޢ�|�xH�z��b�b��WV�϶!�ϸ5�\�.p�^�:�-��G"��¸8huO����ݽ��_|5^y�L��2̍Æ�O�גS)�x�=�ׅ�
%1�9���H!�R�/���;�E���R�����Zv4+)%^I��[ ��w!.�^�hTS����zr �#Q����MO�'hE1)�,��h�a��"�N���נ|�y��!��̃�D�[*���|&<��V)�'�+qBY�<�	Ң� *�����m��tm(F���G�˵�9ƻ���;�ʄ.��ab	�P�2Q!(���УJ�Bd�/>��K�ܙ�<����`%N���D����P>��HW��h%
�4ޑidV��,��P��s+�RO��b<�dĒ��T�s��B�8��"�3�/@QF�%/�\�ˌyң�<�ʣw/^&L	��^�Fi���4�IB��l��D�����wz`$x0h��g��d� �K��w�߇Y!n�{�s/�����Lcۘ/QY�8���l��C���YN�ɔ����I��ć�z��'�3!�H�F�䁂0�lM��tb1��і��$�����/�Qљy�/3"�v}�lďu1�lc/{ e<!�	 ҒGҔ�ZW�2�i�a�d�1*
�Io2_W #�d	#�����P���EJ���3�n։xojz�a1��Wʯ`�>��u0�
E����Y��(����Ң;,�$�(c3�F(�:��nJ�ŵq��;�2-;�}�k������D)�VC��E��tT��|4���;�����cg�����;�d�?����t\��I"1��`��{�	E��ޱ�x� �g'T�,ؼh�*¬6���E>��̨��13B)�ǒ4���,�x��$:����V�y$�{y���b�ȓ�xB�b5NA����֭G�����9��
X�Z�v�`mH�*�v��uecV�F_�<��6��(/������\yp.px��"�[�'�%}61Gމ#�RVZ��San�Il���3ڪҳP��rB�Ny��	z/*��B�)���"X}�{�i|F����*��?��OC\��a��kN�i��Z����wI�["��m�ʅ��ܣ��-ӂ˒�
,H>VCޑ��yG��_��`2��O�#ɜ,	W�,�WN_���e�K2�(h��,ȴ��w��Kty�)�3�mό�Gěa�~h�|��:f���]����:��L�8J�%�{C/�Lҫg�Xț���M+��1%pҥ���ؼ����^�&�n9����sa��rV��Cz�7�L�a޾�9d��h=�@Q$/��'���X���&V�#�1N(���CҤr%����׌<mo=��<��U��W�)OJM����>2X�ד���G�8�;\'}��W/+��
�_W�.3�M��aw��1��A��a�Egh2*K��n�[o��/�ڵ����p@�4ʰLdTP�&^�#c5�K��[�J���xMr�"��,i?�p����i��6@�0^�=�l�K@�$���+\�(���� ]A ��k1�3�x$1Q^� �8=-����-����>��L���"��zY�;�R�e0�b�ظZ�)P%$˴��J�M2I��:�W� ��i�d%V&q���ge�-��λ��Q?�	͋s��3��	vI���Rw� �I"�.Ã��<���k�f��l���q2���q������H�,�|�r��L�C���M82_��5�t��3xM��l�Gpx��`N}X��Yn^G�/I���qR�X�{���|{�'Ú7!�q��\�>��C�2��<J���B>�:浔�����j&�JtJz��J�z���F���1P��骽�`�� �3�#�[��'��;i�׆(/�'�v[��A��dH�>p�劲�4�9i�|�;��^TJ��>G�T��M���Z��#������sg
^|ꫧF;v����mN���.��^�.��*�]& /�AW�Fz�	��J8�3��qh ��n6�2�A�z��BݺxY�!*l������|ʧ*as*�����(9l㋁�{n�3-!�;A����Q<����?m<���s�����ؿ��Ԇ�p�7�N��=��(@��I��c�D�?"@��g���d͎�6i*�k+ϥ�-^��9�� � TP²�Yhy'��ʋH.K �<�^2��ȳ/�S � ˳"C�!o�%����-��Ky�px��o��K�a�H��#>2�dY��sg��/=�Ŀ�x/����j��Oe9�K��5ee9|�w��2H��<��&�����/�����p����歄��6O�����IAj�K�q�^�[��S�
ak�Q�)){���+>-H��z���.�^�*���s������,�{_�"����׾��'e�������}Z�a�+�)%>��m���Oe�s��k3F��� ����`Z��˗yϵp�h��iq[�7��ށ'a�����#�".3��H�ٞ< �"y����.<���x�4^�1�̸wxi��~Id��Z���U�jD�&�6_,�m�O��:)#�L��!إ�ї�QAR��{0��X�:� .��I�B+����v��TRf�X����"�J�//�/{^MV̸č;�s�:j��c`�c����v"�k16:�؈��ڶZ���V�#� |�8�@��j�(�լD�9D��#��y'=+��d�}�����E_�{+����^gZ� h�OT��z`��٨,�'���q'���]���kQ_ۊv���Z�DC_�hiJX�6�#ţ<L��=��~M�ʻP��
�V��U�=J��8���:86e�B#�`-�m9�n�։Z��i�_�I^f�M"������$�|�9�R	Z`���x��`�J�{�����~^�̼�����"�1L�ʔ���/���4p2�xJw�|,�,mD�Y������?��3���h&-� �����'C���v%]�/�;>��ܳ]�W��p��e�	D�ĕ�&���,���Q)w��&���t�~�^���,�kL/
�d�D�:i��-��1�#dqX^2��<�i� Mp~�Y`�:���^sdT���n~��lb*���w���#��|���<O�FXx�V#��x_z���L�����-y�c����oL�,�Ѓ��[�'�y��u-!閘���^��KV��Lq�YN�����wh�`Y���v뗕m�u�+�,�2���ĵiADA2��镼�Q�#\�'�SΉ�r#���X����%=�� ���/�<����K���+��x���d����K�,�h`W�eπ=9G��`g��gB`���608S㕘o��h+N�V�^�8�xt`��PԐ�\Rs�L�9�~��Q�40ƔR���8	���X����A-v��G��'�!l�c�!��3P)C֙�R1��yM��f���1ؖ�H})z��W�z�m��v7��~���o~�F�� ��NA�q6���)�yA��k�ܐ�xG\��B�"`y'�~��x�Ixm?����!*?�y��#�m��
�A>���xQ� ��ãF�>�\�Y�j���e�$2�д\*XZݝ���w X ���2$$��Uщo��M�33������jѾ��u�k���_/��uq�yܔn4�{ɸ��)����E�>����������.:��U�V��G���K����ǵ
��5�\�sޡ�*��PL�Բ��`��wLo���_E��"���X������ǥ��-�΀W�ڼ �)�d�d��N���y����.��z�m�9�G�{���5���mZ�y�Ʉ��M	Y6�hp)t�!��+�6-�#��	ƻ�M:�|��h�ֲ�E�8�k�K����C\2b�0��}��[� ��G��ͳ�����)�gL��h�ٚFx��9Mb�!,���^~�1y6�LZ q�RX�#��Y�D	��[�H��
������F"ȑ?�ۃX��(q�ʇ7�+�&zH�.e@��1�-�U<�$��P�H#�w=���P�}f�`g�'�=L�5A��T��UJ��!��H�(��l��p��D-�ƺ��t79נ˱���}�4c�3::�����4u����F#g�	�S훭J��CCٴ�߭��
�A�+���<�F��ر4'' �xR�5gۣ�R.%����>=&-zM|�N2m?�s҇��5qh�2<�g�A��6�/�����|�N�w�CC<R>f�����X��q�8��ju�X�$�E��m�éFe۸%5A�H�7�lH*24҉��ǰUc�=7U�� ~r�i�X �z�휶�l;	�A�����̹���	q�l�)s��$v��Ѩp�"��6�P��ǒ��M��n�I`�s.��`��H`)�W��\����4�أ�8*^S��=�R+E��{�s/�u�;�W-���3���2!H��4ޓކ>=�ItZ��I��+�KN��jES�-T��ZD�����;7�
Ni����^,��D��L����=�R`ֆ������_<���@j�pe���e[�KfT�%�I�i9�>h*�	w�оBo�V^�(=��k���!���&�,����ɺ��#�{����|�Dã�o猀Jȱ(�9I#�V�k��1�rƥ��_a�6i�lW�Զ㝮�@� ��)ż� ��l'
L�.|����=m�G /g�|Y�X�2-^�FH� C�i5�k���h�T0�R��ߪBx ނ�c��R�@qZ�����b�\e�]�X�İ�c=����>׋�lU���Ge�z��^tw|P�M2��Z���R�ٮ�*B�; _*�t%�' ��⷇��6'��������V�2T��Ii[��jC��{dP哆J%�J����Mv��T%.LŹ�n���f��V�hW���~=�111�k�������h�ԥ��#���'cLMM��H��cg/�&ǲ����o ���{�w#�PD��-�@ȗ�����N�U��7v��M�g[Z��y�|��$\׶�"fR������r|p�];n���7�G�~/w�����1�04�E����kxԶ���$L�8ǂlx]�s���Ax�Z����Ɉsӵ873O-��Y����jL��L��]0fe9r�g56�j |v��b7��.�F�P��������}T�������A5C(N�;5��ȵ�_���@���4�)��`����M�&�/e��<j%����$d�9RF��&Q1g�e��ytpo��E�������Y�1�Q�.�RH�.;�yCX���;�l���I�q��:�e�hO�����X�3�2BxB'��2�R�}�j5�g҅8������QZ�n~v]�oq�Q	�6	��U�I߫S"Wa)�ܧ#a����lS�C��\�3H����.��H9D ��E��(���*y��\�vdF����\2���5  x��I25�M]A�eo".YhCj�������pL�Vcd��OFnƎ{��F'�:P�>�HS���4܆T��.`�5 ģ(J�!L)$�T��j¦(�"<PPz h��7:R�ScC1�A8���4����k����f4�ZQ�����c�9�]�!��1���Q��`��^��#o	�8�R�N��g��U���@�x�d�R6r�f�6�m�@������P�w��㚬&Vkx�8�K���	�|`���n-I3�ïm^�І-��Da���4 Ul�N���71���Q��4�]L���Ӄqe�W�kqvz@�a�tbܩش���Q)�Y�FS716��@�L���kw����0����ͧ�~�v��õ�8��ca~2��Cq�7O�3���F\;<�����Y�͍Ft�����A��M�t���ipg�C�W2a?�{���=<��Z7*1�:�Ņ��o�vWQ>��/_������p�JɀC ����,�Җ!Z��e'��~\[�����D�.H�/�t��U�Ǣ���/.��ň.��SK�qqv,&'FR^� l�A(�"l��u�75��ٕ���;���BR���K�^o��qt�ܥ᷎��|��;��À8
"�匭
y��%���Gk���c#j��2�'+�$A&!(쁞l�,�h&��t��B����B��<ʥe�40��H�'1�����Sp]��E���F$��4��'��Aƶ
J�<8����g�f�Eb�x��8��L�bkmz��3�R���=@�5Z�������WEP�H ��1��J�\��	c[�ސk�j�q=ę�'}!jY�޶�
����Õ8;�E�A� �gFGb��(������q�֛	���I��QFڿ)s���L�Su��slN�� �}�!ɟ��e׏8�xs��şe2�g����SK����d��Ȃ��QBC�=`Z�;��: �Fl�[	��������6�\��=���

�rFSnY"=�p�!iEɭr�j�6A��Bl��b`���˅�87;�p.�UR��p��=�cj�~;���~<Dp��qk�G�w��Q�
�;��iw�� ��~��Rfy$]�X���!iٟwm�%�i��IG{�c�O;4뼏�q]�+��b��
BA|�~3bo7���|g�dd����� %W�^���L�� Z����a���2 :����&׈L����GQA��X�a��(�g��b7^8=�̡t&czt�Q��+-�m���Mׅ����S���fC˹p���w'iirr<>��ĵ7by}3a��Bލ�%]:�>L���b�~[���������B��#�븇���Ą4��R��AJ�O���Φ�F$r���LO���B��ff�����]�"���n��{Q߭Kծ7�ڀ\�8WOP@4���@� ���":0_��L�2����eH܃S���v�tv4>zj,.-��ř83?������cg��O�����k2�%;��911��=�[�l��;{qpx���*�:`��l�Ѝ:ʊ{�������7���QT(<5�sɻ�)�B͠)�V��������zĖ]Q	��|zO��=�����d��J�IR���P�٠ y�Ӧ%�� F/o.�+� �]I�����#��O ��s�6�C\��èmc����v�}fv(.��'��3�Cq~f<&��ٖ���zm��ށ�7��ַ����q\;h��+����Po�
����ڬ$L<���������Q���s���kH#�w���uS�Nt���H<�8/���8O�����H�cs�y�:ځ6�����q#���pŴ?GX�z�
8=�
HF����N� Ht��2�NH(�]��F�2�`vj8���o�</���p����E�8�Y�1<�c��*}wk�/h� �7w���V=��ub��'_������?xԀfa�]F Oj�sl<VNP�Sc`l0榇�=���/�#����0U�֯t
N�֦J�~�U~����������&��j��5�ף�R`��3��R����*�7X�	���S.���g���Ѓ�3����Q@�>ǁ���țRM�3ܚQ;:���a�_�z�l���Ũ\|2vG��@����NH���bfd�#�C�O4�A�A�ȝ@�A8r�8bk��N����bvf �=7�1DG���P04b��	�*�c��}�
)���4���KqC�sW�qA�;by����{�2O>W�qb�p��	��]�!_`r7,�e���w����Ľ���ޣ�x��;C۩tp������r��J)�!�yǆʳpC���ǹkW�4��`k��d��n����q�����"����6��l,�>��mW��ti��V��B84��pL���/���2�^�������'��x���6�uk+ �6��C9
-�&�,Ky�w�p�@ZZ
G%��D���NX���p%���?�#<���}�E�WA � �&���F�FpL�������9���u*�U�h������<��%}����Z8�S8��w�L�g8�e���U0
��<l�̛vM���CD�\<@Xxa��2p۪�I�\!�E�w�x���J�N�3'q��h|���-���1��q�'���	��q0�{;X��{qom3�wHۻq}s;��i���pl@t=#j1#��*���}2y�nCN*��Z�xUҘ{lI���|->��������	����xA[#)A*q��U��m$Mc�`I��s���w�w���I�ڮa���Q�yNQ�	!���u%J����=O'��7�����я����O<�_\��S����@.c�4DF L�b�BۛQ��ǔ9�����͵����.o�[{y`�iE���\���8�X�5�T8C/���!riL�6P#�#��cg��۞��O^���'bnf,�n�@�+��'{TU
��������l��=������a�����1�GRap����F��r����9���r��
���ۺHq=^�ݪ����t�L1�����@�(�ۍ8Y{=����@��K�ڝ����欟���ޤʧL<(�=��t=p�q�]r�Uī�
�\��coS�2]�%��^����Vc�NO� �{�Jy�jb.�i�e�ŗFXE^#�|T:l�*_����1�rC��Ǫ�E�lR��G�d�̛������3��˱8=_�{3~ᵷ�g^��_ی������5��F���y�����1��OB�.=4�ƌ	�|*�Q�s��~j�ь/>؎o<�A@S��*�ypv�gv#��j��&�ZE�3�0�*.*U�4��A��+�!���#/\�={:���E5-Ҹ�e����wwy%n߻�+����+k��pm%r����5��;���ɳ�X弅�SaՏ��ZO���ɉ����31:9�em_� �)�4c��c���7�;�X��&[����yO�O|��!nmxSI�<3/��0���Bb���w��MT�ȗ=8��ݻ6U��N
����J������&O����2ʌLf�D����:�܍��Qt����g��p|�������}�L�x�T�_��Y�udt �Y��Ų�r��9���HL769���82�<���!�F= ҈X�L�Ep&6S�+^S`r>�=����Aso��޳�ŋ��Ǘ���t��t#�?�m�Q��w.��1`������	\�1��~�B<�����1+� F!�u���2��h`s�w<��y���t|�3s��s*��㹴8scxc����$^�;��lr-N��ibj�w49�S>������ZCy��EY�C౧ �f�*����ptujM��c(��_�� �����x�sj~2�'������Z����G���Mr���ӱ05�S�1�7W���6�~^�(��@�c�`vŤ�T�ޣ�@IW���|����X��S�0C�
���pZ?=$Ϙ��]3��Zų�^��1��cdW3Ǽz9f�K��x)��ˉ���(-=ҽ��lv0��{U���/��'���oyl,��A��8�c�v����9)BK2���[�5����,�a���1��֌�v�@���q⁆�|5<2��=�g�CO�J�5���^�]�'Q��N���4��ڏ͓:�)����|I����!��)1�A<���=܉#�<�g��#N��l�|6�U����T�w9�΃g�qY<K�s�V-Rw:H��k'P���xߕ������^8�}�\��ʼ���;X�˛[qwe%�?x++˱�����������[XлX��z/�l���0��Q?֚=�֚=
.��i���R,.-�(3X��ka��u,�F�4B�Odw:�Ҋ�Y����Z�+,��e��p�����Fė����Y�x�Yy���_^J�Y/_-�U&���ڨ^��O!x-,v��I��#w�g�m<�-����O�������_��3�;0Nύ�M�t �A�0xA���S9%�7��ܤՁ~��0V��jvb��X�'H�cS�J%��nA�T���],=㭓�FA��	64>�_��M������}��c�r��j07m)����a��k�s��|�~j�5���f�{��U�d���9���=�'��jsH���t�Ћ�㻟_�gΣt��&�"[;Ie8�䦤vۭ5<*s����ӂ,�������~|���z�6���Zh3aF�3�*�^
A<�?DLL���X������N��s�1;5�pBY�f�4kZ�9�"��0����j�g'���clt<w��4��'m~\'/��,���RE�ؾ�|�m�'�&m���{Ɠ�)Zj���i\��R����G9��ng5�������X��zn2�se�..�Kۙ��خ+m��τ�G��ť�1VD9�yx~��̩���Y��x�����'gQ�x�w�)FbOw��=��Z�Q~�(�����]�(a��l��!�m/�z�8`E=��~�����:M{|d�{��T�5'�&��s�c��=�11���:���@'a`��-�@LY"0��)�QXy<zf(Q�;i҇��2֙��cQ����|je�y<��V��I�� �A��%U������pL󪰴ndq4�����#8���c�8����;����<��Y]߈-<�u<'��vQ6{��'�XZ0��8r����M#SX�A��� �}�#�z���^��l����c�8F��*9�C����umB΀��l`AY(^ŝ�t�ھg��.��x;�-��G^�fy���q��ʵO���o����T8��
��	M/^8��G��R;z��Xg�u�q�"!�]��~q>��ǯ���s�=�b���ESVa��v{l
��\Q���m�FÊG�b��ǉ¨��<WT���xа���z+��'Z�A,�'Ύ��!~���ēgbfz�7��#�c�2��5����+Y��k􀜜� un���Eq��5��0��k�64��r�4���	e�B Fa�IDe]܌g�����C���}縞�	�:�s�,-��(� ������+gD#Z)$�G�]Ng�bfk}�Ҏ���X��k`4YA�G3:&�K����3�.�����w>����q�^�4���j:�J;9���ҏ��m�ݍ�ݡ��\�X'�CF>�1
MZ��!8�Q�S'"���tDK�Cy(��vI>z������^\�vI��Hר,���f�9���4�
	�R�E�p��<61O���o}Ϲ�:xk�jg�7�����r�h)o�WH�ە��*�x*�QY��S܃���H��<�����r҉3.�k!k�s(�1�	�;�t����~��m��A�І��A���_�,��h����ad�V?aPy��(��a�1�i����P�2�5�|���Fb�qή�j��86�������qZ���oq��DQ�Y��ǃ�����tK9�����<ʧ���o��96A	��9�%�TKg�t�v**�Ǐ��$p
����yf6�����w���Xr`bp�ߝ��}�a<x��ۻef�f\/�"���j��6B���&؟�u"T��b�E͕��$�rR�:1A7u�<��$�Q���4�h! ����@<H��T@Z����*�ARq�B��Q��n}� ��"�� ��"1�?���b/޸wZ*cL[�2��t�q����%�děu�V� �������>8�B�Gf׍S0�Ƿ�T��o�~�LL9��L��P ٜԑ�tC�N�S%/o���N��{ �Ң�c&����F��Ʀ�;�2t6$xUL��گ���4� CE4>g�_x�l��^�+���g�i{�Ǔ?�/<
�&�f�\�q�`�Cz����EOD�ѻ�����5������M�.6QNi&H_�9�>T��	�/��|���]�ϞC�;�]�+�p0��7a�-<�M�B4����7���:�)<�4��$NO-�Ř�v8?7���
����<��[I &gƥ!�����@9^O��w>{ޜ�!���1�i(cbMc36�ѝ�z��س��1xxXOxT�
O�����(�9;3�r����f��w��o7\�E�1���yS�\��;��8���u!�^���u	�0�ɉ�<���܎��Q���N�q�Z�; ��Z'&�$�����p��e��f�WQ@�R
�Y��olIGu<����exj%�A��9��X|��OM��Eh�m;k`4�G�)⁌�������!
�R�B�7ʼAM�m/墟������?���{*FG10�GF�x��G�LQP��>��.&u�����¡�Ixj	���4k;�lB�{( x�p0g��9	sw�2o�1'C�����3��\/�:��8��/��?�)��ܝ���r�C|F��h��!n�dL�9��a�أ!a&�O`�-ş��'��O������=8�x:��ݏ;��6]?8N+R�n���;�!˖ N����q^C�l�ܐ3�g�Zď�6�.,�%�$:�ұq���G�ȹ��6��{�����=h!���x[�cwg�W--՛��2�W"�6��=�/���u^𯻜��D����.�f�����ᆲ=�}���#c��@"����N�;�-<�E�Ga����{���ĥ��s�bAOK'�(p�0�������Ql�`8����pv������a��R��n0'�8[qi�T<\~�����V��NiNEĩ��D����A�������O���c�إ�����0"\�w�4`�z.�sǋ2�XG���A� Xy~����-֢Ll/��p��&1N��{�[���%[h]�����I~��������p|Ǔs����^Z�#���Iӓ��p,鈳���M�QM0]K���(p��B�m��PX�m�>�9���J^���ׯߊ(/g%��y%T�k�����J�w��p��O�����
V��]�3V���v��;�͝=���N1������'�6��xpƟ���zӲ����������X{Uu�3�r��0�c6@
4@ʑ1�C��i�X.�[Pڷ�z��d��(3$%}�O�Uh�J�;6vҳt�gm��b��ۡ�C�E�YST����L6��h�.�TA�T�4�৹�8��T���Ϡx���� �ʆ�;��1x�ZC�O�5��:��7�4�|�,=�[E��A!���5���T	)��k�.d<�Q�@9���\�:=9�*�(/GPN���VT��U�r���CA9����Jܯ��� m�4h�a�hP�����G�@s&��	��H$b�������ȿ�>�y܉���0�E� ��TkS�l�|��rO��4)�a���a*��w>}��Il�����ոz�nz<�X���!����i�|�b
d�a����;�Ȟ�S4�](z<|��jxg��\���j}�=���qā���(VJhbx,�Q2��s����G ��`	I� ��J����W���S�@�a�_��x��w��ʡ�J@�0Y��������X�|d��;�4_��y���/}������\�S��[��jG����b$�ُ�����q
!owZvM�x��P:�bw-��|o��\;˱��s{#�)��C���,13m	�<��s{����V�c�W���B����\@�5*�k�N�s����x�S(G��2�Ӌ8�㭓�v�j�F��k:= ���CP��T��΁	j����)g9����z�֞��,�T������ĥsS�>|1>��i�]Ҹ�v���C����]`;ћ�Rg{V��EB�𕊴�i"|z�9a�CG�I����6��9��W9\F��O�U.���d5 @򿞻<��G��f�+�$��v+�Dϱ-�P��}�%|~��µ^���ޏ�T8�5eIs~���vYI;zi'�//�`�`p��ǐ�E?�0J:V	r%���WE�$Asd;q�l��&�4���rĄ����JQ�5;���b����m"����nIY�����ӽm:�?w�E�+�x��(��ŧ��>z*~χ��)*=�i����4%�����
9��h���q��8W��x�0�S��W<���q�r4R4LL�ގJY8�R�ޮ�����\�:1>�2�xH�G�����x>�ggh�����yv�9�{˱�ڍ�k�v��q
]�itEK'��3d�#����	xW0r�~����6P>?}�A�[���F�拆�R�Gdg�`5�B��o���������O~���.��P<�X���۷�������vmcU@�VTK���Tj]���Pz6��ҵ�R�$��f����6?sZ�6�|��㏂
H�@q�y �V�8�Gdwҡ]xA*�����hc��t��
�	�8�)j
�J���lz8Moc��L�
u�ъ�?���w��<���g�z�G����]|���o��ؕ�`�<tE�B85x���x�Sg��F��=��z1ǄC�v�1�QA��P�
wjz��ُ����	�*�&5;pb�9�sj.n޿w�v�u��n��gk�
�PW�C �-�Y���>=���bi�i���L����ƎZ�z;{x�NP >��|�].JV9	�^�UG:��(А��Nk���ll�&�ɑ��Sy�i{��sj��O��w<�?��+q��T���'<w��Ao��G
v�_v-��Wك��"����FG\4��Ө#����:vi�����k|,^�y=����]�Pj�E��P$�cQ3�����{�?�`_�z���\�%o�|l����«��ݙ*�ȇ�T�N]w�Bڍ��kMh��Ux�Ccq���x��;�wr�a�r�����.��9�^D�q�7����$��w���DB*\���0��ʑ|s%8�|��d�M��Uz��y΂��K�G*w��\��!��rXY�
��D|�ǖ⇾�J<vn�� v�f7v�9�m/���\�{��4.�GO����]fz&*��A��Kو띕i�a��2�q��4w�oŻ)�ĸ����Tf�3��҈3SQT�փ�m��*��$rxs{?�a�� ?hC=Yg�}���L]D�m�̛��G
�D���h&���-5=e|��њ���D;��kmxq2��������l|���y|�܎�o݋7�xn�_Nkx|d"&F�P ��A�[�*����PIL�-PN�vJl�Y��
H�m�iE���t�	]�r&��''�p5]��7�I,�q�l4tK��������q�̥��>�c�1Vk�|eѵ� l d�X��a]����� S��C�Ht�x�ݧ�M��^\>��^2.s��|��Xy�c{X�Ma;�`������t�&\��7mj�d�����۲�b/�=����9ꎅ���	�O�&�#�H���R(j	!������Z�;�lڵ��=Ɛ9<ԋ�z�x�(/a³��?��q��D�X�< ���!�#̬/���H�pn2�'`@=ޡ��y����>;�G00�i�UW�����&�C��ä�������9�����ŢT�������cz%8�RT������	�g�]nc������,^ٹF��*5�A�ߘ���Q=LM� HN`^�d�JW@� ���GAY�jo��
��Z�z<{�b\��c�z ��xW�T)�Ί�.CC�J����T�O��e�� ���.1�U�(bZnW�bBA9��.������
��)b@:n�8ՠl�
���g!;2�����NpX!q1��Q-
�(�x�x�a�]��秧�-��vM9U�*ې۾h	*"�c�-�6'�����?�P��S6k��^�\[d���O�����n��x�����O\�={e�<����8��� �}fg�ci�t�M ��k�x$����\��-���B�/,���R,,��9<�م�������٘������@�����2p8F^c�566�)3�nP:�a=X�SJœre儘驩���!��4�vwb��Z�ZY�[��%��{��b<~�B��Eg	ɶ��5F횆gS8��(���g{q�9�ݶ ���ۊ�.�!�����V!�>�qc#�><�?�-��[��}�xlm��[Woĵ���QL�N�,�TխE)��j
5�@!�>��*��5�]iŭ��]���Wc�X]�1��N͆ �����ԭ,�2��x���X)����<���q0��0�4�����k�Y2d���K+Rd�2P�c���ѳ<�u2�։��5F�.6���:�e����	�}���� 7�۴��P"��T��+�66K���2;W������xﳧ�'�)���'�����N�ف��V�΋t��tbw�$�<��	F��d�977�}�*>���9ԏ�177_|㍸�՞]oC���Zԝ��$�;%?}i*~裏�ť�E �*��?j6S)���P'�C��c,G�_oF��&�@�i|@g��Js*\S��7gX�c����+��>��C��Z�.o@�O������K��������;���Mӎ*quW8���u�}��0�0��L<:�==u�8�t��Ӑ�դ�N+i�������@��I�,Ʌ2�(cbf����8{j�*t��/��H������vJ�~�' ��b;^���;'��*G�x3�=�6J���`'��%�6�⁆��n]���BR��VSbٍ�S(�(�#^�&0p$�'^��1�I�!�# 潩���\���F���(��^#���bڐ��a1=��񎆇}��FW�G��r�ɉ���z,~�۞K����j�[ߌu�kpQ*W�\�)�
�6.r΀A�9��!eTz?���s��qV.fOϰ�Qy7Ǽ�F��6��2��+��̞L�s�(��K��;��onm�f}��Fc�7���ݽ�؆.*� U��6rq.���<��G��&nl�����nS�EL�l\�PK{!�m4iC�l��CLv��^��xn:>���x,6�Wcyu3�?܍u�n�S0�,�e��
��V�;�O�Π�����h�IE�>�V�k��I2��C��8a �	y��fHŒ��Fa�$L� ,o*��t��
ʱQ��񘝛��g���3q���8�p:�N]���j��ZP+��-�k��԰!HВ�I�߄q�� ��k�dL��Cn31�'	��F�����P�K��C2]��SXy�����H8��I��m�kq��p�]�����v��}��k�@����0�:��לz�2SO�.g�.�Y"��b;}
��$C�X�0tzJ�c0��h-�g���,!"�K{��o.�s��q����x��`��v�-BZ���_���9\x����)��#��c&������Ź8��� _�S���I,�q��˃�%��kULK�3����1p�7�Vi��@�TV�w֭�7�ŷSƝ:�D��:�Z�I1��-jT�zb����t�^��3�q���S�/b/A��)@�Q���F~*�6M�8:���,Ă�W���v9��\X�!:� �s(�'/�M��xZX�m�WߋǗ�!���������u
��[���X��I|.��sZ��P�I�(-���69íK�}|i1��O��<�5��>�6� �\@�y�$���ͳW�B=T�W3�.���T��t�3g�AO]-����9^*����k�@X��j Z�זQ�z9tn�릟n�c��&�������/���dl�m椕u��#�¹x�|���C��%d���V��y�*Ǹ��枠g4A�|4�W�G��hY9=3��S��Ih�Y��^ em*.�Ɵ�G�P���xy��n ��3~0(�e��'��'S�#�]?5?:�����۟y:�^Z�8E����xs}'��'?�a��e2�����d_F�.J5���s$����sВK��3]g'a�悑���(����1�p�,���{q����V�����6�3�u���Ժh�q�4�=Gc�"йy����D�'�S��͌���l��P*�I�h �gHe����k�2Jj~5>Hv�H�c�PE���y��sg�1��E�r���X\�q�c����8i�c�2�:��	܀\@61V�%1g�'��xϒ�ĺ�<�x�'PDv��^��2J��liO�3���g���J�ֆ�}.e���9�Og�xfb�H��X��S����)��!�#�#�:��Z��Ba+�fc�4?c �&`���TOp��]��Ϗb	�Y6�sAw]����o)1������8	B˙p*��:�D�;`k߳�Rr݉�M�f~f*�Kve(0���B{c(�!hibj����נ��NL��N���A�@�\���X0��8�uB%�4���D&��bA���JZ�Y���y��8	f��a�v
obvn:�����4�"���CH��3��TTS�k��c-(����9?ǀ�_� ���m�p[*�����j��8�q\smn��4J�B�f���S�'b�)����E��G��s�x*�Q��Qxlj\K�كS�'����>���1zn>��D���`p���\�c0�a�4N��c�nr3M�5.�i$�eG=�o�64�#!�y���h���+�Z`�,_�G� ���2Ьm<{j���8%��ݷ���!������3�rM����on���v���Ӱ]<u*g�CWʯqھL��3AI�wv�M�L��kiXkt�L��kڝ��f��*��7I~�G���� ?�t��* �����-I��:�!�ȚӦ�5�-���j��ˎ��a�8���S��>��x����[���A����'ď��Ff������l.�,����l�H��D� #����o�c�w��+�+����]�'�D� x����7�.���f� l`x22��"B7p8-��J�s�j� �M��i�a�Z�P��9��R��LO�`>zG}o'q"=gt��bm���Q�!���-�B�5=��q��3��3��SO=��9�>AC���<@��E��<�}>LY����Rt%r�Cl�h�����SB�A%�߼��|=�c|yV�
�xx��`>�m{�I�����RϧE�"�\,6�F��48�!j0Qt�P9��Խ�Q<����8FO����]1��9���R�*�yr\�r%������4
�P��q��k���LP�Sh�`w��U��Y���TC��������ذ�v��4��p|�YX�
����dd-Ca�n�����B���ʮP�]/4����A�P�v�R�^��ދ���VO��QOΙ�*����!\��u���')\���X(&q�+ٞ�36���!5��tp�6����xpIz���)�s���A���D ��S�ws�d�"�Pк��&h��h�iʟ�7g0
�7�}�`I�敳�=vg:yB�i=�$�ҼT�ލ���m�}>>���c����!t�R��fכB�{�/ӥK�	�($��k�S1�8$�|�8�o�L����T�\:놁�B��%qBz��qn�o�_�?�
�>�Dc0q	�T�_��L��~b �<9�|υ�鸺��vrwwg��Ah�={>�kk�E����3�v�I�emN��S���4��w���3�7���TNT@��|�l��u���.�R�1D�2A�*�qb1%��9���N��3�r+�=��]�a��3g�c�_�S�0p�*~�@RJ���$N��\K(%�s9����i$ ����^5"�΢����S�g��?�����D�ݻ����u<� ���T*"x �k�.�]a�Tl	�cw�8�LdÄZS����˙������ѽT	���ʀ���Ԋ�?�/5�)���Ǫd�DN�=8;�ۆ:s�l�����������+��r�\l���ې�k���޿���䞐*ȶq˹4 W<�#�Wlx���K�adZ�{)Kj�^��0�G�M&����5����8��>ha����Ȁ��O��y9p�L�vo���/�}��������tl��\ঐ��*�t�p������b�bL���U���8>���G�
��ۀ2���B0�@�	��X����a���	�ӂ��d�q�(��;,l�܎9�o��h*�mC�E�i5dr9�YگTE����<����LR�3�'�� �w�yd}0��h�4�e��$T���ý��{Vz:9ze*n�ya���t����h.7ihri��x�`�uL�o��LQ��8i���f&Gc�PumH�:8������s ����v�9m����z2r�(�#��{�ڧai�t2���> �x���2���8�ͨ�T2��>��:��Tr�Ƶ?���܋����+8�,�i����.w��Z�>��^�^.m5Y�g����.�`tŽ���zCv).���(`e�c����z98-c?�єP�J僜��`O��q
/H�85U�C��%�!���1O�eǴ��᭬vv�md�ť��HFp�ܜ�m]x-�����}�1P��g���sQ;M�9�Q��B�>���N�<�k~>�L��*DK��ܲ�� 蚮=����4��.��O�ſ��'���%��[����7���*Ќ����՜����Xk ��3Z�*�9ǁv��g"��na�
Lw���������<S��Lo��`L�@[�+	NK,�$&���S�>��Π�/_����c��������A�Q�ǰ@�|J7��`�^^E�[�;G*��xY�����L�r,4��q�o
��'�+���+�=��2�u����^�K)2�lF�7��� ����R�����b��x>i�c�a��
@�
���Kr�L�)u-�)�-������A�Ա� !�\tKza"e)���oif2Awf]�������������-�T����4�2-�{`V	�]1T��K�W�rz9�ݪ���a�q*�'�B{+9�((��j5�\q����V�lr�Q�0G`g�UɈò����OOp���_�Qq(��8<�� �W!�3{���ۋ:��vz9�!�)�T�pO�
�����,��z���|{m;��H��[�?d�;�5@\�?_�6� ��Μ5�)�a<���X�ى�k�Q?@p�}2äO��la#�RV�vlwE�g�ZvG�&ԍ�bG�W�6v��=�_��^"�\(^�wJ��P��=G�Ļ��3�l:�R^�+��nœ�#�it0.^��?}#���۱�u��vz��/��Sg��+{��Ёc��e��;�0�{<U�P���i*'�\�� G�����(�C�}������}I�ԇ�9����&����ޕ��a{�7�obt���I��4;�_\��s��D��䷬l�^$��A�&_�5c2J>� �R#�W��!?s�$k	N1%�vy1~�x�����8�h+nܼ��=�o|����S��Ǡ�׮> �PgULN;�m�RQY�PI8�,�#J#��ȴ\'�� ���;Zۦ�)�~���L����6�֨�Aan�9r"�P�@�N�����3q���x!�'�[�X�v����(�J�
�k֙�7����׋"��;��ɀYFa4_+w2e�^��g��ܮ j�ˣ4z�)g��q��T�wp�q����^�G=�\1�P��>;8��x'�Y^~�3k�c�Y�B E��1���g�+�S�Ǎ��%i�zHO����)/�JjɄv�VJY�>q��E�NQ��%dw(*,zc*�|�Ixpfo����m�S����x��K�0�	"W�I�Ⅎs����!u$�Yr��v1��	�������\�H
��%����}�}�h���=ګn�� �[s����n���{��{��*ij'�^�ye�i����n�x�._��&�Nl���4}�y�A�"ЅАx��z���j� �����z��{�֭��+�����������w=:�{4�B��mS����o+��!��AI�Bn�/G�j�l^�T��=�\sίq	�|�k��F��VpW~H���o��=Diü7�������5j�IV]��ڵ]�C�n�Y���S#��{Π|.G<�]ݎ��}�h\:{C�LL�N嬰!�;��4�<�7ƶt�t��c�����ql�^#e�2�g��B��_di�-"p���I���Z�
��;�O�^�N����D���ɱ�����7��|��b,M��π|�Ds�Q|s�h'~"Γ��G��3�k�4ٯ�iy�u�����o�!�����_��SX;���v���w�wr����٘����I,>HP�X�޷[��6]M�Drz!LL��PDj���Yj Y/�<2zQ��l��G�u*]MpK���#�*��]�9��VX�����Vg����v&Փ( ���n��e��|$v�AW� I��2�/���{�(�KW���5��·w��ޗt+��zedzʗ�SA��uI��C��`:8R��]R>�ᠽ��kO��~l2����3 �n����J(�*������y�&�٭D�2��Q#��WW7� 8!�������B���ݍ���y�LktK{��Z�h�j��ܔ_���e�4g�)�J��!M��W��N&q�Y_�w۹��,�m��z�R��xp����?�nu���G(l:��BEa���F��{�9|*;w\p��>���W*ܶ�a��<��
:��b<�C�ƣz3"�v�Ls{�����]
���<������>Dx��R��f7k�co�Oe�R��h�~� %	M�'����b��`�lm'��#���^,s���ٗߌ_���q����p/*�%�^��U���4.�k-=�E��xO~!�픊!�O�g�N_Ҿ�K��{�����l�E�}�e�Ҩ�[�9F83�]?h�.���O/*>p��=��Y�xv*>�¹�Ihv[{~;����s����{Y5j7tayz9.�H(=E	��FB�٦ұ�z
���F�xd�]�N�w����e�n�"Oʮ=��,�eޜ�uO��-����m^���8�{p��=/\�gg'�6N�ǐ����}��l�1����l�v	J-[4VN��P-i���;��l������3�6��յ���G1g<MM���L��q3Qvw�X(r����Z��g��ZY"�2��^E��W�;Σ��n�]p�tE���M�.�-������~��;��������w�X\9%N/-�@s#���O׻��u0!�"�C�#G�8d�υw{e���оWP��]K���l;�zя��~ƗȒ/��y%Hy�ҘD�}*>�2iT �V����]���F'�wr��y����Ew���	ܵ �0�[���d��[���^��G`b	o#�˚
��S���}���xD�QK��$����qq��`ͯ�+��}۾߲ ������������23�����߮���+�9B�l���B���_�#�?9z:k��qw�`M�u�A���.ₗ�����^�S�5����C�v��]�nwg/�vvh���^<�ݨS��vSif�F�����[�}��q,�La=#@`\wsX�:��;���pIf��I���Fۯ7��q��V�צG�@A�w�2��7v�����]=�ŭv�tU�榁���b�C�`���;kkk�Z�reWm���
�=X���
J~�v��Z~@�@���pcd;������,�&���22	�����Ē/-9�}��7����E��/Fw�u�mh	�/���kb�4�	xp&���c>H�����t��u�`JѓCq������K153��zn;D}�>���r��2h��B7���/)�JWf�I%�|�Y϶�� Wy�H��|��ƌa��B'�d�2^�P�(]we��CV*#�2D�����s��`?�W����L\�g&��Xb��67�G�x�}S���(�\��u�L)!Ȭ������x����.�Q����Z�:\݉v�4jD����t�D��ȁ_<�`�*+���"ǳ�E����u��4mV�����Uo&\O�J��Ά*��xOn�[��e�l�����/�P������飋sSq���p}Sc��E�k�;�u0U�T���9�}ƃw����f!ކ��3���^���hC>��6���{eP��T0���e�����1�x��(��v�.�Ǯ�b��Q�~OA�ٜ�0�(���������ڊ=�޽������ߋ�m�H�����0���������.����*�CX�>gP����1ܸ��v��<�O_��﯁�1&��Ĝ���	�=r�	���� �B��b??���E���G�S�N7�wod��sۢ�qW�^�V�����Њ��y��Vp	�4���A?ت�͇�L��OM�-��0�{j�K����6�	}�R���mlmn���v*P�o�n7��x]���bqv2���ih~
�8�/߸s;^Y]I��
5��z��Ж.���׶�q{y7��s
��i4�-(��{��o^��ׯ�蓶��O<���A�H�k������py%�ܽ���ƻ��1���"벼��E4�N�Pt��T��Z�.���m����LHJW�x���.����kh��I������/�5wc�����O�U�B��w�89��>m��RT����R��
8�<X�127�}���Ee�5��4�l��s��ĩ�yv-F1ƩO�ZR��p,u���~�}S6��i8�)��]h=�C�.n�*[�_L	�2�1Wy!'^��T<�����\�"e��8ͫ�����_0j/�d�0�(��NF�� _(�zB�.�G␠���,�vp�˫�Э>ʤ���x^Bh��p����܅y�i��y� ���~�?5�3�&�h4�����Q�W�T���V�*���&�"�2��d�࠙�:�X���hq�}�,�v�:�,���b�BL����ZE�VE4�I������<473O>�17{*F� ��V>�
f<A�8n���;`ڱ
�;d��S@��d�~����!���w`)���{�E�FR�薚>)�(0-贚,�@풠=�x��#o��!�P*�3���䠍����j+�\9�m��zH�z�(w��{sx <n�F��Xw���������[�iQ�I��=�!��z|��x���h�-L�*�R�����0�B������V�`Qw����
�i�k+�����haՈwWb=4�111s�d�N��@���V�57=uK�v����5���O�Q8�;��rZ(F�OP<�����;�hסS�3����'��ݭ���Zq�ߎW��Ϊ럤e=�at����Q.L��&�����<K���Q��Ċ���n�Í8���[���܏C��
.����l��mm�+wWI���@�>��1��K�&�gl���=����5���h�i����阙�̙j[[(e<��x��m<X�����������	
�cok3����<ܧ�:(�I�L
���V�YY�[��q��ns
�K;C?�T>v�AӴ�
���1J�S�MƊ~��a#���A���X�ʖ�MUe&W S��/Gu�#Qy&N�p�Q|�MV������d��ǝ��Lb���<�N�F���Dgz(.>6�T,-Υ�:&�E��3q��bNU�^��&�p{�ʍƞư�#*U$��;��tf��)�~�_�A�^G�rDf��x���.��I9.UP&�-�vθ�u� }�=\��x#�m���Aw��ʯŬ2���c�	�_N�&�]�;�q���pf���Ȧ|��*��;fPp�����t�h$���puw�y3ӓ133K���*�ҟ�����;A�ŝ��Y2�0�ة�I_��ng* ]GJI�}��Z��ޏ����.��dJ�x
.��` �/�M���0s��1���{np�z�A��*����7����/�]`(���81���k�,��w���M�/��EpiuUR�1D.�x& ��Q���q�ފ�w���^�h`[�;xx���"(T�X�K�q�♸ta)��(��@ߋ���؀T6H�՚&+����f�`����-�݇qms5j��8t	��U�\�����B�m��r3~��:��>t�0w�a�mb�CKՑ�����x�x�g�cz
�8�|��Wc��v�M<�@��!�a��+d����?i�b�yW77��e��2��P'��f;0~��w��+�xm
�:8���]�r����v�e����Ѣ��ic1Vc�?35~��Am������p7:(����8�4�xp{����nMt�����7���{8݃A�60�ၥq�yX-�rDA�O�����8޾|x���S�(x
8+(��r�/�4|�Z��J����������[�¸C��I����񒅉�������{H�ц����'�c�M	�E�1A�
�Я��ʧiT�.���������l���ǹ��F��2H���&/Ge��Q;�!���ѪN����cP�mK�%[z!Aԑ��lW�qg�O�cx�~�BOv��%���1.���ſ�~(�D��m1����
N�;��zP T�uv�!y�,�D�~n%�ĕ��:2��	�l�`���g�w�w���2��P��l����s0oO"{mZ,+~��(�(��5��C�����@�b��Ugt��a1�[ɣ ��r.��V*Os6	�`�5���`a~!�ck#Q�Ȫ"Ĵ�Q" Y��vrJ%��WD���GzN4D/�G
���q�-��1��*��2g��T�T>"�
�P�޹��k�6����LNt��*��_Ϧ� �����1�G)-�%b=�#�$L�s�%QT-,rK�+�"3�;/)�:�����y�+Ӷ3���$>�;玽���S�N��[�����(<�]�Z����7���373������g�K��ܙ��Cػ�}�1�gtzƵWU�Q,�Q�Ȳ�QG�n�4�惵���kqz|xA��T��awg-���S��ۍ�ڵ����߉{�W���wrrT,H4� uGO����'�/���D	Yo�M�u ��ctOx������)�NV��x�w�QTZ죔��Pô��ꐝ]�̏j�!<�xh���_�����v.`v�aO����4��?�F�X��xlc��.
j�6�F#`#�H?D�ZX��dm�] �+^�y/�t�~lP��W�ϼ6?��b���v2bzOZ�K��cy�?wm=n�(�x���ql?
�/MM���L,p�B�8���T9��pO�Q\Fچ|�S�:!gl���nn�[7��7��`/gWNcq�����4�o���Zhڣ��޽����M�M�c(�2�%��p�>� NƢ5���y2��_����h���|H'�(��csZ�Sq���si�i�����9�q�8�(�S_���E��,y��1ó8�6L���M�S�x&�{�35y��]uT^���#��*����?���8V�9�R�{jv!������X��4�m��ib�w)�xUp l����N��hC\��哏]�),b���Tp��q�s��Sgs���}�M!�c.0]N/qd�+�<~bd'�Q>�S&��4��rΆ��)S�i(�DI���Zo<��Q�"�[,�I�����1�����y���[&*R�<��+#'cXn?�C�P��}�A�z��%3?�%=MX!�+I���e�5Z̊�ܿ.��A�t�dG����8�Ռ/|u9���۱�U�Gmh"Ƨ�z���/�Ve���m��:��'tv1N/Πx�b�|G�Q��B�O�n���+k���ߌ��]������TT�	!����?
�JL+��E�~�?���������Q��ӚBz��,=fg7N ����d�^pϴ�8��@��D@�P1ZI?���n� �<^�S���������-�$�&]~T!�eG(3� }���T>
��nܸw?�����k˱���C�hZ�aL9~6<�SS1��Gy*��F����%}���h�5�M���[G�X�܎k���so�MY�Q۞�
�Og\̀w�:�W5�EJAԿ;A�Q\�}͇͸vc/^�������pЙ��n\OlLOo��;g�u���E�v�� ��C7N�pwl[y��5?��U|����ҵ[����F[/��L��(C�T|aVd�[5��B�b�s�s^�C}Uz$8����9��;�5��xoM�F������G<��-����UhN�y��uE�:�v��<wr�JX#ͩ�I�	�;��L������J�����)=!�5^y��q.�m��1���(x����Ͽ7�8=;.�Ɛ���LR T� �# �߻!&I��������j���2i���p|ཧ�e�մ�],&����z
Cf�b�����m�;"�~�qK]͜n�"�(�)#�������5=���ۀ���Pl*�0<jB��OT��:�n!2�5?�L��%�8�8� ԟ��e?&��{@2Ż�O/�G'�?��_ԋ����_�£0f�V_?>˰] &]k�t�����U�ڦ�	I�������b�V��+_^������^�� ��S
�?!g2��5��|�R�⇰��s�G!�W���mB'��ݵ��K7�'_�[�����k���u��>�a��}Ua����;ԡ�׎��\���׮�KW�ю�T~��������sT�~7�}�f����@�� 2g�h�JHf��a��X�� �_�z/^�{����(�9F��O�d;� ��������y���j�/|c#~�3oǫ��^z�k�n*�%�_�]�lK4�Jݱ'�Wu�Z9�жk:9 Og����V��֝�;_�F|��h�!��a5�Ih�
g|<(�	��uy_��Y1ύ�XGA��k�o,ǚ+����D8��(�]�M�n�i�uE* Ⱥ�O��r<:��	̯���յu���w��;��o\�7�nE��\(�.^���A}<�LY7$� /�_z�I��9i�	R�U~K��G�|�q%���v�qzrGN��B^T�%��Ơ-��k�X�E����У��ymn����1ע���:��
��[��'��c��'���&˴BV`�x����v{ACD�Fi�|��K�J�����߉�Gw8~�07}5r����x�!�ǐY����/�t�{�����:+X*'#8ޓ��41.�{�`���퐛;�6`v�4:7mw��9����u������ؐOE�SGP@�-�p����]q*��z`T��#��L������"�-���O�WT"�S�iQ�N�w�9��t��kAI�.(�"�g=x߉��<J�-�ѫW���p��W�g#x�Ÿ���_�/��^z���.њ�
\���v!�����8̇��:�y����g�t=n�ߌ������ĭcgR鑠 de���U8n�C[!��>�xN.�S�'�zl��M�������~#6� ��x�߰ۆ����Ҵ�D� ۩ॐ�h7X%��~��7����y��:=��~'nx
����g��F�y�t~3�v�O_�)�*(y��77�����ϼr+���V���}�e�I�xL��F"y(�Jk7���&�
�
�W[񳯮ŏ�n|��;�`�z�'�2)o{8Obf��qiܺ5�;8�=0m�=p���76�+W���|���4��ѝ��ök�Ǣ���s���Q��:�D��xB��uQn+��浃��/ߍ_�⭸y�!Ɓ;\C
e�u.���q��
�����h�p��A� vP�7��㳯�
�o�k�6���D�k#(��������,����@i���J�д�K��?:�yN�LTZF��.��aU�D%F�B[m4��Y7�u�M��l��&'eY����J�f\�U^���[��ȏ��3��f�x�%<�#��
����r����k�ɮ5��������{�74����/�Q�|�éq� <�Q뫱8��I�C�:@�qy��D g㬝�m���#���r����x��v�v"��������v9�eh�����_�q#�w7�瞎ť3Q�>O�]ׁ2�
Ʊ����A������u�F��8Ka�DwQ�	4�;FTV�|R@��o<�E�)�{�� ��p���\�����5�7�?��B���apUk�^���� @�k�㛠�g�Xp��ض�0{o˖�{�z��12q����Ķ/L ��g�Ѫ��eс`r���d�E�M,�kG���N����ىQW٨�6P�)���rU>eFv�P8(�/������v\[ތ����7~��x��Qt7��x��)^���<WQ۽7N~��Eu8��#=<��N>Dq�q�-m./�b%vr��OA+DF���Bw��I'��`s���g��S#h�~+[qgy+^~�a�,��o���Cp�⩶ti� ��]+��2UF� h(''�]z�ծ������g�:�	�@?�x�p|�tx��R~7�?sK����ճnuZ���Z��
_�ʫw��//��8i�k���P,
��TdN�?�"lmx`r'��%?x����J�p}g'��b�9�d�]�ѝ��\T����0{�C7�[�}��7����+�w_������#�=6G���>��\@h�u��ђ/JF
�.��Gd���yj;r٣䒮�H������7�ʥ���=�P�ʤ��!_�O����7׽�7�P�Yob�Q�,mp4.��o}�Ÿp�L���]�?�.,��̨^� T�e���ØRt��Gi�7<���o����7���sd���^�wn��٥-/_{+�>t�5�g���o�G@��8���j�3G~�~�ϣ|`���^��nn��.�
֚�0.Bᅋ�o}�rL�h4ԅ�ߺs'F9�#����h��,Z�b���(ʇ3,A ��y%V�X���}���5g����GRq�{�d�~������yda��}�~vC<X�o�vƘF�\�ቱ�YE6i��,�:X[���IR	�#���82��)J��&Ӂ�<K��gʤb�CK<��<L�c�=
���d.˗��r&\�h��r�5膱]a�G;׷v��1��v֖=C�Tf�|u�Wn=B�~�_%���a�;�>\�_�f����Z�ܯ݈ի(�{X���t��,�d��إ]���X�]YN�� ��_��cq�|k�8�n�Ǚ���2�{��ĺ�P> ���=ʩ�ni�����.|\��wV��(��{�n�|c+[ ��:��0`�a�#����Qa�U>z�*���8>⬽�n��=>l�`\�=���!r��K<� T�("�~�>\�@�;:���m�v����7no��y�f���a���ҀQ��gF�sz"f�C=3ਂ��Q�~�&���]���~+��Vk�۫�q������,��&��e�MGE�R��� ڸ���������x��������K�h���(G�E-�x.O�e�DwoMza�� 9~�*q�n�n��P�H�~�G����������2;N�0������P�h3�n7����=�-� ���-��T������~t��$�9��߷ ϝ��{ƭk9�pqq)�z��J��@���V���Ł��P�A;fj�}�S�%��������[�¯߾~��E^{��kq}u?ַH��(�� 倖r'���˽��qv��X������A���F�~k7�*���uQqe<��O>�Xz��H��d޼u;F��s/����׬�{L�v9��w{͛}���ɠw� ]/7Fٽ3���2�� ��ݻ&���w�G����w�y�^l�o �������U���S194c�Sѱ��1�U� )�:è���";1ρp�F��-�h!D�Ty�4O��CYg#Z��D��T%ѥ��2����SH�Vf#��dH����9�|dW������~�������*¶�k~j�{�յogA������E�Ž����g��V��_y3^��W�~�2v�|��ѝC�,BW~��ǩǀ�Q�p
���ER� L��b7���5�[q��~|����ǂ'�3������ݵZ� ���n�_Y������ڊ��6��W��O|�z��K���f�v\"0C&���d�0|�x��6sN{
.�J�H�ٲ��#�ܵ��׊�G���^��c��������:x<�̓���|em#nP�7������Z|��Xc�6uk�Cޭ���9�[� r;�A�mRC ����D.3V c�x��e�ZPE����㸍��_84
�!�� � ��m�6���rܸ�_�����j|��X{Onܵ��t��.�� �{�Jɕ��F�ÿ�Y�q���X�~��E-�ڵ:�;]�X�;�4k}��H��(_/m�~cr����
�E�{D��˵���<$�/�[�fӭ��j����?tOg�܎�+�ɐ�gc�'����"Wx���{��?SD?�s�o9������?���}�bew#��(�4�5�o���i������d�ȉ�^�Lh�29�����S;�����zϧ�W�4+-���b��O<gȰ�� ����B�$.]�BÏ��	����c��Q1�B��B[�&�H`�3�}��j��*�Q��7�U��d��M/"/��f�oݻ+a�[w��՛�Xq��X��L�iJ�֬��E0�v~���=RN�`��؃˾�����Ē�(�w�/9�����<ػ/]W\Y6��9��xoC(N[�R�7sѤ�*5��~� �~o?nll�X��ˮ��م��ְ�[�h��o�lŗ߾?����?�o���Q8m�?q.!�Ɯ���F����,�6���
��I�V���.+&-9}8vObc�$��_z��;���U O���_������.�r5^{5~��{�v;~�++q��h��`�ǈ���`��u�C�!�aL:v�88�HPh���)���V��Ҕ�"�Q���v�Ykė����>^�I��}���͸��o����޾?��v|���x��X�Z=������|�Ľ�mK�)�aω��$�WC�KQ���l�\ͯ0�#j�O�݊�A;���㵷��+x�������1Js0v��k6s��_}9~���l�՗��V%Z��k����{��P<�� T�W~��)���-�9�6��(��N�l��Z��yJ^�m���&��Eّ|!� WԿ&��R{���F��T��R/C�L��C���&nrj ���b\<3��b��s��q��BN2I�\
ο���w]���7�A��7=�����aG�܍{w����8���g|��Պ�=����V��Q�y�3���.�n����;5���#?�M,���X��nm�;�~��)�T�����Sq	!�@����wnb��+W��Ht�	Ys�Y�`o~/Ʋ�im�rd4o�
� �T6D����?��w�����cey5��{ׯ݋����N,���H��m��'�d�d-s�GQ>ԕ�H�Z_v
$ed���ګ�^T��)H"e>+���~��O��댗aL�(M�>��:a'JS8��Fi�a�C���R�WQ���;�xp���~1}s7y��#�Q;��ݸ��_����7������D�o�u�t�Tĵ,s��9���ƳC��5<�"L�؍��F,������]�{/9�"�uy،�����k���oߏ�������1���v�'�v'��߽/��J�|�$����4�C����-7p
��<9V���[�k@�C�'��UE_���!��e�v;Q_m�������~|i�0�nW��F|��a�2���/����qxoo{e(���xsd���1��GaN��:c���'7�eI�r_L�ly�Q��J�/kx5�#?A�+li��~%������xY�z���u���6��a|�����~���쓧���f0>���|�s�v_$ ce����S�Ht)�Eg�C^C�+�Џ�.)�a-��&�'[���<S�S�	ڨ�g���i3yNނ�z��q%xM��iƽ ��(�
?`�W��F식��O|���������A.��˻��3c�]�,t�]/��������^����8�0���q9�n�1R�Iw��OkR�Qq.rI���ԭ�`LMf{�T�&��B+�fƂd���E��{�d�Ȅ:�?�q�L��/�x�h��)�	iy�5o���2
�)�)��>��c=(�����������t׍TZ�K)ӕ�ś Y\��zœ5$ޮ6�|�=����ZP�c6qL�q�D��8�)o9�Aʘ���6�"���w����"}n1��8��:�̹�>�]��v�v%T�(����ø�Q��u�8���܈�����?���}.��G��o����{��F�G�� ��� ��6�<�j��������1$��d?\����9�`�<����6^�����
���Q��۝�|����_ٍ?����č�w��k�?��Jle�,��Ht�ɵK{�s�k�՚��3�lK��pۂ't�:�/5�\;[ʎ.�:Z[9WX�#��̍+�;���o'�W�Nݸ��ko���5��!/7�xL�[s�2.���O�ɹ	pI��t����n�d���@��w�E�����M��(�g��s<N�����<I�{H}v��<��~��z%6׻����x��@�z���q�vC(
���7��D)��%�\\��ѹ�uF1h��cMM�OA�䝊�k�Q=�-9� q��WjI���:˔�Eb���&�]�I�J|w�s��e5��!�'�ݺ&�S(�����#'ϐ�]j��u^�ؗ��=��p<8~�|�/���l���I�ʗ{y��z@C'�?w2�v�N�~R�I+�q$���lK�g��:�zH�K4���������9_���+{�����ٲ�4/ x���ٙ�Ά��~w�{�v%_S���7*�B��,����PQ�ZWx���.���9�j$jx꙰��I�\[�a�[Q�o2H*1�{����?Li�O	��>JR%gw�2��d�|ɶ0��{��]�ٵ�
�sû!�i���mL��Ϯ�����F	���B	�:]��*Jkoe�ى����}7����^݋{o5c�f-���� �c�ha0r��A
j�0O]M��-����O�D9{Y�k}�3���*R	�o���2J<0:vE[��0�\WY��]�d��Zf-�x%����M��덁��i�K5
��*�v0���$�3�q!�evY㖑�11��I�ݔb3�c�k��O�+`s]Q� &4��MO�2
��lT�h�U�|�C֥�a�O�~���� % �3�7�SՎ�U#����\��� 7��* N�C��XoE����Sʮ���FōG38��Y��'��8C{O���-,"?���Y���1�;�^�G H��mHD�����;#�(T����DI�m�,K��6i�&�eɅ��^���g������3?�>/f�,����YYZ65����;�������L����|�Tĳ��{8��(nܹQ@9f	η�vb��n�lUA|vW��k�8/y6^�A2x.�6���HHܨA ����^"4Sd~~������N:������hp�~�)����Lz���F��?���I�q����>�G`���Va�A�P$�+��FV]}�h
R_�W9�A�W���H��{��5rQ\F�#�|�J�� ��n)���2S���\�ЭE�XG��i�#�����[=X��|Rqd|��&�`�NG{v���0��u�A,x7�@�I�i�GzG���x���ּ�Ga8][�Vq+�Zpg�,6q�*g�J�R���fY����/u��\����0��C�rLcf0&��it���;~�Iē�(	�N|�c�dg����b�8��B��:���\&���M�������9z��S�Hp������u��Õ�G!���[��ٗ j�K7��V�� �,�~
E4���@-��O�k]��Nχ*�@����B���1X=�]�w�s�����h_8��%��Gw�����u&�� Hƺ��M� �����)��1��)ܓYp|�� ���A���p��8�A�u�R�'7n��v~���Q'���{b�����ŵt�]rz��g;�T�x�E�di�����6�ے��
�5����Y?��J:�P�Mww�p7�wcnj:���Yx%�~lS�?ᇟ�p�h����n|��ø�=�i��c�έu��׿�t�G�*�9����i$�8 �b)j�������e��_��F��f�U�~@�M�l�~T�@۴I���ov��}�/��q���6���2���Bgى0�˃:Z?��3��P�ߣ	��3�b*q��r����S�La��D��q�!�i{H�u�����P`* ���yI�[唣P��� ax����L��vA�,4B��Q==m<�j*��٩�3�fV�1�G������P�:0������4� @)w�L�:������QpgZ p�� ��H�ϗ<��R���hn���k� �Y�pq��p��y:���$i���vqFޖ}�\`0�bU��(����޷���6�4�]�H���դ�*�4� ����8q 2�s�!��HLN���(�(Ȝ nspG�q ��C��yψr5��u�����٦���]��p��b �\��#p�w��֭w��8���~�=�=��=�ݯ��NEgq�ұ�o�<�0��}E�A���|�31�!�ը�)Z�#��%֦��8�S����AI��l�z��/ݩ��AZ�u�qL���4{~K	�h�����W�'d�=����K����d���P&��h�LcrO&�DJ�&��S�alWG�?t�=������~n-6�Bж_��Țw{� 3�'���t����NLB�n>�����sud���#I���7x&��#��%�k��Skm��z\}�'p��u�Z΂�������mOA��csg-��R^+�^8k�1����e;g3h�!ZW��a��F�H/��	�-ktF�c9����߈{�o��7��7oa����;#Nc��z����T,Y@�C��E�Q��G�;����H�`'��+��*Z�NwT_�S���ɣ<��*5��r"L�/6��@h�XN�i�.w�N"��d0�%w=8iF�� ��<��f1�,��T^�1�+$]5�2��t6�8B�A�&zj����� FPj�Dz?</8(�GϹ���pl����;J&��9��K�5��G�͍���Ÿ|q!��K� ��:�M��"����	nd*�N�@���]�+�X�è����/�M�9��"L��l���8��b!��6c`�3[�N�OD��h��!|熐�s1�v|(���"���k�j��=�#ܝ16�����=:�)#�1��Q����b��S%�5"��b��L�?>�L����X8������Hϣ8P�Ҡ��t��e)~� ?x�/��m� �U+�T��ef��Ǩޮ�Z[�SO��{����<1O�%=��\<����O\����bowx<����q������J��,���ݳ�T�~LK�wg�i���f�g�OT�*�ݸ<|���y&�>��I��]̹���� x��b�~v:��|*bs������Q���Qa�D���[W㭫7b����w����n�����x��i��x��=��Y)gD(7x�13�<j4��/�_��7⧾x+w�((���������|2����\\y�y��7��|�KXl��=���X�>����u}$C�v��vc	��֢�i�!��4J�#(1��w�Z�w�;��(}�ĭ�'�����_��g���k��_)^���hξ'��"<}v1P>m���2D-]K��p&�����ߤ`�U׼�q�����R����= S=T����ٚJ�64�&rq5��h�`Q�f��d�pp��F�#0&�P��!�����C�W�D�e4�Atg�;��qtj6��ӈ�=�K��'8cx;�Vt��F��e��O78&ӂY)�۴���ߛq�r=w�uG�0J���� �x�8u�Ui�FAZ�
_�^��j,��,��Q%�]�ݑXD��"\��ڈ_~�a��͈�6��ֈ�'����b�xou/��oE�ٝ��E�	ʟ��y��T���ww��c&t�F!��_F���F����r���=�0���C�뉞��QQ4������:^��t�f|��~�����O���ѱ��/_����]sC�?y!�M�����8��z�l|���x���7V�o|�v������0�~X@+i�37�/�ǿ����ϟ��q�W@��5\vo���s�o���oū��S/prf,>��K����� �|����џ-޼�R�݆2��P'�_�����w�����������Ǉ.�ğ�}�ŷ\��Q��ޮK˕�>�=B��~��I��Ͻ��Ft��>;�4ȩ{f�sm �
��>9��1�Gji�k�<�}v���8?���g2)ʮ���_duAp��{;�y�nT�!�]�R�}��3�~��N�{[q<4�}��x��<E`��Ļy���a�=�R��{7vᯭoŏ��/�Ko��Wczl*n�l�����j-6v���d�W�4�V�qZ�g��zJx���g�|��>e�ݯ�ی7�e?~�0m�^S�z;�M��3��ⓧi��X~VausY6�K
�4�l@�Jn�QR?E�>�xt�@�H�(�~�o���x$��!yX��:�~���x���q��J��ֵ�E�צ���TL!�G�P���7�(�U�ßb��x����^gwJ��;oI_,1�G��{G��24����[���),��_<}R�WO��t����?>��������F`5�H�E���&�۟=��{N��z�T��N�~��������l�>6����@,���P-���9�^������w1����x��ɇ�����L���]��������^��S�q=�!���b9� ��q�Y�ٲ	`R�����u�w�3-F�����c}O����d|��/��x��0����^��<y9>�����w����sg�
��.y]�w�^����B���#��/���X�<؍�{�ݒ9��X��&�O��|��x���cl|,�ղ��W=Q��9I+e &�������z�����&�~�<僋'/�O���x!>�����S���Sq	/�ŧ�����XA~�`+���?�/�����/^�{w;�oث /��0���Ŀ��~�S(�����e<��n߉����M�fjtN��c�O�����?L�<1]�%���h���n����!$\�Թ����wc���(��G�Ŀ���q�ҏ6���av�����Cg��h#�wi>�/�v>�zzlv/�o�?|a&~�wQ���A��f��/�;��Q�gf��3g����p��פ��m�����e�����Z��������\%=i��2�����ףn��{
]/{������%
�8�j����:4R����g�'���s�s�=<up���W�o��zX�GGOqy�`y���˱���16�_^�݋{;��m��1H�(��<R:�u-��8V��40�v{�O}�/~� ���w�0vףq�di�0,4�8�n#�w}�>�A��~~"�&�Ȥ�n,�����XZ\?wm��� ��.�~�[�V�"�:k�[��ŻS�V��[�R��X�/Ӝ۱��o��J�{p?�-ߍ���?��g��X���12�����z#9�<��vٻ!}�aSE���}�S����A�v���g49jnz4�A�/}�3��/�mwu*8»���2dP<��,Mƿ��+�����'^x<ֺ�����캚G)� 
�_�$�G/�w=��re6^Ċ}����O-�w������x��*�m-����X�Q��w=���|���d|��������O�p1>�����{Q}:��+k�y�N-�o���4*���1xW�h������bW����{<N/��s�1>2�>4��Cqej4NOWc�����D�l6���^L�w|�l���}��K1�^[ۍ[7ע�$S�K��Q��ޟ����Ɯ]^ߏk7c}g��Ɠ��r,�>B�]C�L����d̏c�n~@qp�����IL h����q<�w7ZGq��F�ꝇ�6�������|,.�V��DL �~�kw���Cy1zy.��C��o���ųԫY;��㈟������v�{�g����Kow~$�<3?��+����̘�3/�S��=8��S�_A��f���]`�`�,����{�Ww������]�/m��}��H�������Ӗo���Ǉ/��o�<��A�� �?�.�S}`��ᄂ'�����b|z'��CTr .k��C�T��^~�7��\�'�<e[d?�ͧ�3��Qg���G}���$���3�� +ۍ�v�ނ���O�sg��Փ8h����L�@?}`����=��z&.i������W�_{���{Y�ɱ����qoy�`H�~F?�Фk�q�����H�X���
����|���~w+j=��2 9�Z��'�w85=5�.�K��G{����F;�'Fczv
7F���tȏ\�:��ed�vy��=~�T��������C=@L����o��۷b�`7�߾�;G(�Kqؚ�\�鉨b�tX���,��o^�%]����~�ę���y���oqv���=N���4.c��3���w���C�x��v�L���i`�Lt���8?������R���xey?fO�ǿ�OƟ����E���&�Aol�S���3���%<�x}��Z/���⻮��G�	(n�}/�>�j�Y=�1�k!h�۱O����z�o�#��L�	�혒�Kn~�����)���bvr>�����_����|&��_�|���?��Wbcs��(!�������Z�����}s+果�O>}.���x�`?^���Yً8S��_��C�Ƿ�E�K��J����իw�aW�`��t4(�p�qoį�l���W�>����LF��+q+�������W���|c-��o�_Zގf�|.�xBO-N@.���06����͈���}��_�����/9�|5�s�O��ڍ�y����Svc�H��32Kg��O�R|�GNǬp�n1T>������x��N\����$<6FsL�oo5��Q=�wq:�wa:����=9?�x.o�ًʛu��,ų���Oόd7�Q<_z�=7�k�憵?um7~��^���g�Ǐ}�A��7��,��ubx j��O��]�[�_���jĈ;u` ۝#�>d�j���r��|�I���s/(h3/hj�y��w+�w��Hp|/�Վ·Ҳ#�| ���/��E�l�MP��ى������S�+��NGAY�vB(��k��]�{;>��/�Ts�V��7��q��mH�5i��T>Z�6ͻ�����<����7�ϫ�_�ėP>_W��O�U,o�*��Z�n�!vFF�����/���׊ݽ=4�Q�n����Q7�zK�mS�nvW�8�\��C)A�{�֥�������k-gZ���=��7�o�|;��6ce}3^{�N������1��mzz&*��5��<$R��y�M��&p��
�������UƤ�6��9�������x��X�=�_yu%�%�]?�b�DF���OM�w?9��O5!�7���+�{���g�_���x�� _>��/�܉��n|��J�~� �w��8��=��ÓF���Al`���s��/�B|��F�@�o��oݍ��S_���Wc��F��A�m跐����֎���q��7�W�3�hN�,�Zh��ű�tE�i=sn>��z_BH��U��{9>�߈���ۯk�������X�p�T���O�����U���<������8=;냃q]ki/�||��Ғ{��f|�k7�o܍��c0k��mn��j����@k(�{��݊���S�'1R�=��ǯ���'~%~������0^���o�������X������p\�˛�`���t���^8�?�����{ӊ�N�@?���9`�`$�NzQq��I�ѝzf6��\���S����?���������ތ���r�Ool��VVb�w�`8:��m��+o���q;>|e&>x~�(Z*==qvn:VA��J��V�P8����x~6�����_]9�/�؉�b�|��D��.�/��0~�o��~y5n��7��ů��M��{���:у����"�6QVZ"�㴠����J;H;^(���]��^~t�n�^���o���xy%_:y�����* (�1�}�̹�x��aCŝ�g!6C��e�����IR:�ҹ��ߋ�~�K�����E�/M�G�}�x=�ñ�;��^��-='��WR���mFd�lx��-D�2>FI���ZZ��D/�pSX~�m���Zo����ǽ�ne^����D4��x���u�fT���(l ư:`<F�i�����u����I�������2ͷO�����{��^f�:�s;V�@q&�F��&SX6]�Lg��ʵ�8�`Z�r��D���K�30P��{�Ȟ�C6�����1Tx(@wt�;Ȗ�O����CY�L�� ƀy��n������}�cq��yVc��G����g~���w~�����W�O�������?o߹�V��z�ӣqa~$���3��fs��><��������o����ף�����_���O���_�L\�v������q �
��2�cH�ĐO���!qH�HnM�Vg�묫nLO��7�1t��x���z� v�^������a��xq���Ҍ�>��K���f���J7Z�m�����������[?�t|�sO��/����~|��X����Ӝr-��$|�ثV���S��8����=��w���Q#6��X=iŽ�h����mD���� �WP�(���UG���ފ�n�d��(�?�G_��}{|��4��X~��n�������T,�[�%��a��P��,h�u�y}zu/��/]��ݏ�������\�k?����|;��_�z�[��K�#?�j|���q�"��m�؜>O)1J��Z��o���+�\}@yZ�z��CX�'MbҤ�o�����D�_9��^0
�?x�A|a�,�6�:j�v����w=��Uk���P�<�?���#�TL�-��qjt��]u�l.d������a(��9�����G,׽��{hch|4��V��W��W���7����!�6������7�b�z���2k�mx��U�ҏ=�[}�k_���]G��1��@�x�1�����'�GіBܕ\��Ч��5��y�[G����!ގYg`���0PWkz� ~��v���݌v�r�Ҧ�bvj��q����}�v4�0��IBn#�6!��P������7���|�f�]��wbcc-޿��{�����_{��<����i9�u���N�R+Nx)��������J��!���{�<e&ι^���y<w�� .�$�p}�����'\bi��ݮ2�� �9X��c&:��}w��X�������x󗖣�U,ͷ6��k���Y���co�����������/�+q��?���8?��C�4N�ڍz�|�8��K�Qy;�kG��/oğ��.������o�v|��ר�x 0�D�g��5J\�IE�8+�@=0��Ve;����>�%�uz�f4[���9����*h��gB��)W�o�7>���_~;>��h��yl2����l�k���8a)6PJ�W��oߊ���Qٮg��b��0��;�SN���jô/���i�Q��Pt��v�M�)��tF��]gp9��w��1pk7�w�J�o�՝NN5��ㅑ�����J|��Χף���Z3�ʏ}:^��WP^��O��Iu�+�|o�!�؜0��|���D�����XԞ�C�~�?����W������K�s�(�BG�qÅ�m����8������'�se"{5T��YIHJ�>��0�����P'~�\��6\%�d�.��=�͚��uygn�����TM JR����
�.MU���qJt	p\jp�gP��W�~���=J	ri�"
w���X�'"fߣ�QV5'X\ߏ/���٤nx�ׯ_��+�i0�Z{���"�
m[_�)�ҫ��K��.C>����z,�wc�p,�p��\���>xP/3H���hm��KYe��JʲM�6��	֛+B%� ��־��H���l�=��|s-^y��bA_��Ν��� ?�W���]�M�n2
�I%'�� ��QBJ"*���E���<4|������(����|��wz׏�����p/<�kk����wooō�;���p�$8��c,V����y�7YG��lTⲜ^��|����H��J�^m�֬�S��m/p�6�u5E����ڱ���F�d�ݤIs����n�,<�:��$4qx�e{�]i��G�n��FaN�bww;��A�����?����k�c�q3�41�5|�[w�=ރ�P\�G�HRj{���^|����K����v�STy*!:ȍD�<�����9�}1���̽.��^�/��@W�ż_�D �a�q���:�iƐX���9I�w�q��x�G��׷㗮n���Q����3��.���e�m[��a����xsz9w��=9'̀D$ER��E٤$Z֒��l"�,yI�E��R�,�4��%AI@ �1y��s�{�/���9��������T����{׮��_��]����E�|�����`�l����/@���MF�sbվ��� �8W���^58V�i1�G�tR빇G2�;+p��X����cxy-���w�׿�F�Ó��@)N���W��zm���������1���(��n L�u���i�ǰ��C�-}
��1� [����ٙ8�g��G��C��_�+?s*�?{,�>��O-��b%��hOvi���~@���6�ez��G����8����W%�7M��K'zx��#	����D	%�/����z��t=h�����;xP.���-�e[�b=C�q�Ȓ����s�z�R����(�d9��sEh*�]<C�?���x�s�Jr�<S�G��1<�l���Չ�71Xᗗ�oD�t�'��7�!�¨=�j�0�#�~�g����D����_p���~��w����nC3/��r��ګ����^(�`Z~�q���wH�H��T-���-p���<>y�!�\��;�h�%�!�rZ(<0�!�2Q.�t��0�tsM�/�}��a������Iw���8�\�b����fܼ~~9��[�;�����������w�_\�o']t��Ї�Շ&=��?te�7mF�����bc�Flܹ�;�qs�~����8����^�:���@���,�ݳZ�92�ﭖ{"� �2��88�Xz2vB~�wE�|H��_��3u�Fq6�R(���S��s�8�����[��4Ӄ��<V�z�|)~���rQ���}�w:�_Ɗ�9YM��
���� FwPL����{�-`���Cfx_#��{�� ��R�UB�m�D �*Pj6$�H>�0��,h#�/��[r��Q�KcuOE�1�ŅJL��Q�s_rsxg�3U�љm���n�%Z�{�ظގ�e���m#��i�Y��:�W����~�ո���c�*�!�*"���	W)�o�&�.-UX�S���d�����r��WF:,-��
+%�n�\��"^���+���wi�x�=(�Tz?xi=~�׿k�)a�WV�ν�x�^ě���S���u'&6�Q8=` 瀆���V+Nc����=_��|8~��W|�_zW\���7�������W�O�ӟ\�Z}s��!4�:}�ýAlt��.�l���ǧ�;�cst+8f?e�@��kq|�u�[��Ĥ�����X�"}xZ�C�`E���]<�צ+��<��;c�Ɇ�3���"����A#j��S����Cȡ��!�U��l����C��2�O���X?���K�x?�W����om�׾/�k���t��ģ}��x����ǰQ&�?�� ��:=ȭ�;���;��f�����=� ��x���⫯ĭ;�c{��;CL;��ҹy^�N�a�o4E[J��2���<|�]Am��9�
��/rɵ��y
��{ �B���\<zv!J#? 6A�������lƏ�����F�f��L��7oǏ^{=�ܾ��v���`� @�X��ҭ	X���A	��
M`%N����d���#[\z]��Nd��H����xn�m,λ����y��fܼ��ڽ��D*���l~�s�
0y9�+`*:��q �|��t!CA�~�|w�G��"��B���C.���E7]�읚��/wi�b�O��~�mROcB�<�z�� �S�q���a�kX�6ww����t=WI!a@����{Қ/vGЀ�'�]rI�*���|#��X�S*%����ڴїL+�՛�Ҵ8=dWe�2z4ޡ��������5�f�.N�f�i���w<������:�s��ѝyzL����B)�QWo��w/���>��E����a|���q��m�3^#-=Q���G�G�hV�L�6?�7D��5������^�~��v	�}����8�өJ�[Xׯõ����V;}:�.���߼��PV�AWc�b ���-��[�1z�C�
�W�9	ݪ�ܥ{�֌w���Y�+u��q��gf'�g^��YM���)��{(�?xm-�|};�f������:x�d~�X�.Oh��_���R`՗s�����$�/�ҷ��39G���*t���q�#iT8α��]E$f�{��u���1}�����׾i/�����}s����R���R�o��@��6�3����cȈ�z�����^���������h��sq�1�ۛ���+�����vs,7¢�tхߺ��;H����y�?v2�O�:�%����x'��GuN�2��/�/��r�ݽ�[��;m������8��Pq��G�a�1��G�֥2:���\E]����p����C:��v���j��#'��O����Z������������Ͽ�Vܾ~�"��ر՜X=��p���^��w��U��V�i��]��G���#k���  `R���B  �C�	'���?q�w�ѥ �p3�޹���7����q����-�����鸼��.�~����v\n� C��,<y�>綸vw�g�Q�?��w��<(�xX0�ù?[�EP��A7M�S�����o��v+���@Zn�B'ٔ2��t�D���צ���ɨ�(�X�c|��7���5ϯ�
S�l6�6��|)G$A�`�M�Sp��*-KI�C����mdh_ĥৼ��uQ}\W����?��>'�w���������4�:���[{���������Q��[��K��:��Z�0p�04f1��m�>�c/<JJ�š�n�^���L_$��d��~T�RL:Y	x���4���v��8:��0n� P�u��Ѡr����"��h�>jUt3e��I���(��s+�$mӲύH[�l�Ó����D|�3��eS��ܜba�F�Q�_��9E��q{?�����7�(�3<�ȹ��~z:N��@�Ig�(��A/��`�&�w����%}�r�:�o�ݒ�{�9pycO�Uc�O���T�qԁ ��QzUB. "�C��7����x�]:�@��d] �S�Q�q9�Pʏ^�Z�r5&'�uѿS�����K:��W���w���q��_�/]ُ��D�v1�����x�7�ʍ�/�;��0��pғPYu*P����A��qɓ?~\1���ؔM�{��>��y!޼�<\߈�a+7,8�u�x���n)6�\\�1�Q8t�x����zX���1>&�I�=}\�����G�
A��.���.D@GA(CGL���}������۱v����>�s�Xh�������?�Q��������eJw�-Ț��8bq����M2��分�&d�>D����x�ǏG�� �R����Zܺu#�ܼ7�ߍ[�����w㕷n���[Y�ٱ�Q�5�S���*
�A��"CG}��o���>7!��Q*t�+�`K �:I?���<�+�7~PΧ�G�s��:ݍz��C��<��D�ܡ؉Ow�Bq\�O�}s~:�u����n�2��(_���|c?���nv��L!y��T�C��
IekVՌ��u��=�!�C�9׀��Iq���Y��_~�)�m�0f��\������q�E
hqn�ˋ3�X-œX���GN����|:~��S���'�����_����C��H}u�Όr?���oF��=�Bh����B�gg�S��蹕Xp�4�W&�'�>�~�bT^�!e�J��h\fz�l.�,�T��hW��[���D�NO��*�o��	���#��hR��i�8}�P�?}������@��kΞ|r5��g�2{��c�l�u�t
����Ѽ���k�sp�ֽ�������ߎ��+W�˯ޏ;�*��]n�:����!T/��$���N|��Z���wbWo���B��gf2V\e')ыPmB��h�z.���3P~j[e���9dc��z~�!��Y��䙇��R�8I��q�c�l!1Аԕã��)�yrЌZ{#*�������R���Aāêɗ�D �֭K��$�	�ɽ�P@��Y`�S  ._kƗ��WnbPL䢓�jm�ƕ7ߎ�QBw��ajG0Ȃ��x�s.$#�<���V�W4G�>Ӡ�&�=,����ݵ�����Ǜo�V�y�x�|�s<�^'v[�X?���.�ء�d��U��{_���,q������o|�g��5�T�7ltB�W�1U)G<[C���U~�҆����G�F/���~+����A�lF�>�R�9~<V`8G���ߎ^x9���jt�v��H��#���"l?��sE� �QBZ�R��.e�I$���(Nq��S������Y�3nݹ��z;.���_�_����̎�|T@е8 �Z(H����W�9�\�0'0�,WFȀ���h}:�L\�y��	��A�B^��r�m)���u�D���� WapK����U��L=��l��f����f��.���<�g���s?�q�s���`��� *D�x=5Z���<�"�g���&�1�����)�s���&�2B�ŝ10�S��eN�:�ơ\�!���+���McDcC¦�ݴ�ዐ�>���^�x�t���M���U��}��ݫ����׶b��6�q��b��L,?��^���48��>���;<���>���c1un>-Q_�U����f�
����O�'(�hO}��C�����<�B�A�L���j�Ǫ�X����>O�^�x��Q�3d��?s���?�\T��{cP��̑���0���=W��Y�&�8Sq�2^�/O�ᷭ^���/ǿ��_��o}=�������o
�RhOѹ�ގ��o0�vZ���W7�Gw�?2P%�_p8_��ɝ�i+=	�5p���r�Z�X��(%H�n���N�;���.P2���k	D���(�������?4�i�%W�F�`+�[W�t�[1y��Qk�Ť�C�a���e�?�L���'��s�0hzB����\� 3�H�����n|�7���2���3�zgȟ���sC�����kW�~��u��/�������:���!n<�PqM;����Z���Ǘ���xᥗ��o�������nvۣ��⹳٠�k(G��-d�l=�(��B���a
��SWʴ�ʚ��5��eaw�ȎKO�-s�a���|��$g6p�sҝ^.���;q��0���܌���Wc�~KrW��W���Ṛ�v���^�W^{16��E��ݥ��ߡIƧ`KK��tz���MA�;((�&����bwg3v�ec}3nݻ���D�܋�q+^y� ����y�B��ȓ����+��|7@OG#��QXk2ٌz����N�&��iWՠ�
\�f���v^6V&8Rd(,���61»9�q8�0z��+���J���|"�.��+3Q���}r>>�H-f�6X2�|;��hå�j����0����y�M�~V �p& #���}��b!�"��Tc�����cb�6��G�	h �/�n�9D������Tz�n$霏�F*~��#q��C�̕T��_�kŭ�^�;��(V���'{�a|��~���Zv�C@ʯ6���W�/|�B|���p5���Ɨ^_�o�r?v� ��X�y�R|�#�������8�T(Vi�ps�å�c�HƁ8��+hUU�I�y��0䀛a�偒�܋�y��R=>zv)~���ܴ�w�.�������ާ1�?��j�՟}o���1�>��c(��E�xj���31��,�4�&�ٺ>S���cbz%�|�Q��>��(n��)�%�l�F�7[��@����z1�ݍ��~?��܎��� )���H���(L���V)��E�d7���,Fs�ॗ'b���&148��{���洒uR���$9�cZ�����x�1�"oz(����W�{�eh����weF�``g���"�?�����g�O=����T�A'1 N�����)��3����qkc�#C��75:��M�͛7��^�?~�x����sx�;#hlùG2���_r�L?9�����^mW��_A�|��ߊ��|=�޼7Q<-��"��0m����D�ڪ!��).���Y���S��Cv��0X�ѿ���%Gl�y��`��V�b��b�@Q�4J��{d��c�3XVu�gC*w+�y_�ҋ��kW�+?��k��j���c�q��\,OOE�݊�߾��q�ʕ�\_���f�li��.�%�?h�CO�T��������"�ωl�Ɋ�<����<���C�lnlĭ�����7��k���⥷�p�8�� ��1�d��ע>=�����(�P`�t�ꆳCX���/H�QG N Q��D�
H/�H		hZ�v��Mp�@%�q" {�NM�� �n\Ǒ}dy*��O�����1����yf1~����k�=�@�RN�r_���we#����W{b�e9�*Gxk��b�G�2�K1��bT�c��� ���d��p���B�ly��а��3�(C�>'��6H��\
mӳE�覓ٽi��xR�@#�y�������G�������/�0�ۚ32*��h���`�W���+�3���'��O={<�߿��ſ�w����G���D�g���GV�w�����\	XЦ?�-��f�%G��!2����<�&����U#O:j �:�C��5\.�c-�g�X�'P@�,7�ͯ}�Z|��f��W_�L҂�e��>r6>�S���S������G�a0�Nc8��"\�\���8������ӏF|�\L|�|L_�=�z�CZӸ��Z�R��@P��r��v��gp{'���n����x3�9;��"�ҕO�-�`�5??}�����}�L4>���,Ň�/��:�E��2���5)��=�/���P��i��t�x�4$�=֦c|A�Vm����[8�1�JQ�xC�6���f���Wpa��d�M�U\�����,��h8�"]��W�z��7n�+�{�m�|�WX_�f+�76��/�~��ދ/��z+���Td���v�X;� ��(�A)�v��6v(g�u�_����Ǘ	/��r�_[��������������Rl4'��~%.ߟ��u��Ȏ@~h�>����ԡaB%t�W,KHg>(l��_<��sq	�1�����_�hv���6��k[X�H9���ӥx��j�z����u�!n�`�¤/5�l΁���zk�[;T{�.���U`�9�O��!.��G�lom���n�\=gC J�*��v���-V��� 0Hj�+�'q�Od�lT�},�����V��:��{������U��s3��z���hq���V���B4*o��aS ��e��5���#x
!��B1������
���VE�/��[�t��ǲ
�L�S�KH�� �`z"�Z��i��ا�j=�s����ss�/��d<sqQ<��K�����z����qX�}��,ʑ��[��߄!�2�l��Ђ�(�O}�t|����j��9���sKq~�R��U��w��X������e �G��s3���J|���V��7|סӁ�$@�X��5�����Ԯ�;��h-�o��������byu!޾׉���k�{�:̻?��Y ���ա9?|�����O�Ճnt�oǪ��؉���,�E9M,�o������Ǜ_�;��T�qfi:.P��o(����ڋ5?�ʼ�;2Hu
9��~����]a$�e,�'��ǥǢ֨��[��G/]�ݵ����p��
�Qm!�˳��|����.��csqH��q�0����x�^���T���B_�Έ�U,G��Gk[1t�e��P��ڠ����~�:7'��b	C�����3�<>K(��Ǘ�=���?��P���f�����x�͍xhe.���*e��ū���b���[�N�4jѡ�gW��ᕆ"C����xm�߻�O���fc��, �?U���F�>�O|�d| ���S���E�D%*����-�o~����݈�Mq�t�Nb�	n����f8�7НV69$m�,=�F_�^��c0w<z�ɭ��B��9��c���SA��(�>��3��C龆����p"ޟFh����F;6�Ѡ.��(=�%C1t�(y������B�!����"��e�
��%�B�r���8���Ho�"W��N�޿o_�?x�x��������6�;�nw0�w�nC�(F�s�Տ7����Y���,��xd�ļù��	wp)�:g�T���]�����e�<�k�c�����O�����/n7���[���͍���ǣӓ��ç�3�/�ވ�.��ɽ6��!VQ��~�V��?���x�^����Z%w��V;� G��M�-5��V����X��v�znJ���1���XB"����bś�@C@v�2�M�� �A���:��Z�� �nx������_��߄��^���wp�!<<�	5{#�Ҙ����|LLa�C`��o玴��3����okC�\����2E�>�g#�/&2)����A����V���wηP��搄�R� �k��nX]5��*D������*
�a�A�p� �_߸_��[�Eh_���Y����`��ե
Jk:�*��/�c�\-�N������_}�|�k?����ǟ��Ņxic?�NO,��yS�J?�}�D��:(��J�>�5��b������O2>�ާP^�ho5㭵���,����h郺��h�㠄� z�z���Z����w�ԧ��;��G_{-n�v�����o�Ǘ���k*NNW�
d�3����s~�X���/�6A��ڊ��[ߏ���K1��c�܉B�"mY�,������^�Cg(q���#sѯ
%M�bN�E�?�\���tܼ�_}����K�a`�(�jҏ�,96?�s��C����[���F����-�9����J4���[(�^��_�p9�N�F�:�ߟqY�;ʟ��h�'P��9�?y�T��㯼�t�Y����sr��A�����o�j�6�]-�O>y
e^�+76�_}1n�z�.�ق��PZO.���&��D/�ڏo�������Bݱ������K��O?���c���ŧ.���] 0�Vg2~���������aLІzq�����-�M�\�fԗs��������)y�e�=޾k���V��8��p�����%ɫ:�y�y �Sɨ�'[��֝e@��֘��⢬\�b��Q��k�Z���Lç69@P�w����*���wbsm3�ܹ7��ĝ�͸G���9���[��h�0����c��7�ދ�w�oxP������x<����k��ى.�z�����a���� ڹ�q}���3(D<9�$<�+#�ە��-p�ovm)�Ls�ƪ���b%��$�."�,g�O����ү��t�;�ү���d4�F�=~�X�@�?������@���%��TF(���wWFX�~���^+m:�FV��\�1�Uր��3��e᪖~�����۷c&��ݡ�]s��rMwA�?�&J���m���f�;t�iv�Qb۱��|�F�����9�C|�T\�X��:�ݸ�^����t��`D�������������t
߲���+������)t
<8'��$��+C���G�|��$I�t�����/\���-E��K��� ��K}_��8�Q5�D�ܤ�\~�4S�U�i����UM<�76�������_z#6�ئr�\��q��K+՘����q���sx9/��?y&~���������x,�����ӌ\�?��oS��v�>��ש�D}�x�x��G����C�^��~�\|䩓���U��+_{1��k�r�t����و�\���#� f�ߢv'ǖW���i=�o�o}�Ja�%����;{�n���	�;�mA��7���=�O^:�>X�����|�x�f
S� ���}:���|fi��\�|9�F�z�t}���R+����L9���7�n��޾M��}���������r����8�H=��{��Q������-���D��uz�ԋ:���@?�r'��w_���wq_)��-�}����^\]ߎ�[��R���*p2��;��rj��Ȁ*0����޸������k�iF%�}�d��K��n_�|'��͗���{cEW�)��N��{nq.�PH���;(��9��腅X�E�H��ur��#F�,���w/������_��{�`*����~�Ȳ���s��_,�!M�����������i�i��oB�>(� _�Rqq��<�ؐFc�)�ɋD�8Yr�on�r�e�q�z��}��xB� ��OA#e�uH��'�9<�|�6��W!���{w��շ��շ�������o�Gs�֭���k����A��&i�����]�������E�m�N��r׉�[U�t���n���T�٭�����N;�5���m���L�}6Z��wh��<�Q}Ե�|^��<�l$��`���|�k�?����XT.1�4G8� ����*Rl&(F��G ���3 ����iMƕ]��X��sAC��U�:^P�3�FL�k:`(�W����^�o����d{+�D�67bog+Z�{�:؏���Vr>�Q��(+V�N�@(f����h��i�y�㭛w�7��W~t=n�6���j�X���b8W���z�. ������Tz=P����T��-x 	�p��h�T@`�F��Fg�:�뽢ϰr]�[���IҺ�$I��H�`�	���W�o�bx�K��^�3jB̷!NW�,��b������ލ�����{(��W`f�J���\��^�"_��E:h �)�cK5,v�r-:ш��j�\��"���[q�N1*�hceۈ�i�	*v����Q�_��ՙ8{r�w�[�^���~k�����S��Qp����4i�
�%�=�o���
"��u�\<�oa���Q%��O�o��-��s�5	^�bH�tg7.Ä��F��(B���y���n��Mp�p.-���t�7�Zݸ����s?n�ۈ�}�hU�Y!�d��yQ���?zB��>�&n�����ְ�ɜ�E@�UU��
�G;���[�z%���=���C�9�M�-��&|0Ө�շ���ft_݉����8�-��u��[��u��vF9a��s��wsk��l���z�}��_����������5+}��tvq6.`��G��ƽx�{�b����2�E)�;��Md�|���d�:��W/o����2�pf.�1f��}�w _���ۡ�mڴ���۝����Z������_�l�/H�Q���\��+����C����/���5p��4@�t�0u��ks��б�{�ǿ<�)<+��c�/�(�!�8qL��;�����&�/LB�.��l��rg
���%S
���A��2B歭����:��nl��B�ܻ/=���?x9�ѻ��ƽ����ڈ>e8�����; �x:w�'�x�qc�mb����"��)a���Ӿ���F����7@�=�f����T��!�0i�Y�'����쪓�?�=�����f�Dx�E�������>�w���|�Xϯ=��8���Q(�D��wׇ]��)T2��+�Sqf��]��{.�ę3�F�!��)���� �t�#9�ۦkg;*t�4�]���x#7�ԛ�!/�',�q�����sЊ[xE�a�˯���n��0hi	�-���ը��ٹ�����+�@6�
�� ��߉��r�S�G�n)Z��Ɠ���w����b�ʷb�܎�G���OG��m���NM"`i�/�z+ts^��ݓU��q�sq+v�܈����"�=��U��Q��N5�O?y<~�}��=�a�Vl;~��7�7��f\��Q)��p,��%���n,��|��d\<>����HR]��V��c	��o7~��o�"�q��jlM4h'F�4r���g�}��5f�C��b��|}#~�+?����BtH�9˻��jd_BU�Q~�4�-��*
!q �]n�u�~���0�r/�����1#�?���/���cv*NXn��s�db��ۻo��9	t��--k	��f�B�<��DpXF����
�e��\�Ri:�輙x�u�E��++9����m<v����|r��oT'��N�2�����x�����&�ڀ��@����O��SO��M<�?���6��Ҕ^s����(�ƁF���T.T�����އOҎr.�ҘFw�� ^�ޏ׮��[��s���9�|nq1�57��W_�h���m�v�\�M��ǖ"�9�]<Mz����y� �����r���ep�K�����6��b|�~+ׁ�>�Z�J�V��]+?X6��O�4ڤݜ��<�R��*����Wa������p�A�q�{h�T1=�yTx>�d��^�>�}Υ%y���<t Q8�I����Ȏ{�;��	8�1�Z�X���'J��8£��-c<��=�����MHC*}�L��A�����BNj�k��_��P���'� o��zt�M��)�f��үF�)v4��]�a*�?��3r�G��4�8�k%䖻YMg��ǣώP��z!��7�Y���s�3���8u2J��h��ͭ��_y#~���!�V���S�|w��"�6�ՍV� �&�:��L��:0�nc	�1а�_*�r�E�17@�D|�хx��<t]�r���j�kO�� ���tZ�kW��|#����.�*A'�L'��j����:W��!��"�~�~��U������Awp�i�h��#�������rd���);�꜋�#z�v�{;F�_��d#�/�/�GY��� =�bY������}9N�c���F���q0��8�"�D�0�ʠ�u3cG�3��S��Uu��s�n�\��m?��9q��1<v!�倂��B�?^�<���u��W����^��d���
Ŋ�,�����������{/-ű�
i���Ľ��x�[�����Gq��Xz�JL<q6v��
5��:�<����� w0�~s7�X�w7������koG��$ʉ:�,馰��x`�S8��\`~VH{ ��Bq'�&L$���ښwj(u�����á h�Q�|��7�b]8�'�����# ��G\���p������K�]U����i�ؿ\���FŤ%�w���MiFKZ�Ǐ)�"b��i�p���Ry��{�I/���������\��-�`*�&P�+3q��|�/��h�Jc���C>���[>�����>��4x�Z�#<����Q���_	��D��-gi �_��X^(�@U�.$�@-���[x�й�)���"4�8�qn5x��F�6�8�Og�B�D%�=�/VOg�ܙ��uC�(!}C��B�]�	ЯÏ)',A��\(�Ш���w��#��	�=���H���q~��W�LBw��RL8-����!?A%�x��C{9۔���pz$_!�Չ(����mhmuc/&�M�!�TJ�tr2N�����h�@	9ʁ�Q3�ݼ�rdj/����y��=tO�I�*��&1�����q8Y��'c�=k��	��E_���~��)��̀��< ��T\Y�8��P��3���b����*�PlZi*�>�d&���/��1�N���h���B�|�g}�������z66���o른�G�\��Ce����txM?Dӎ Lli`�Ұ��R�Y���g���	\z~�c��@U+���ĠY4�|ģ�@p�V�J�/1���u��I�\��ŕ��;���{�q��F����v+��XO�i,[>�g�u<�w�XD���Fyv�8)N������>���E��?�(V��>�sρ�Y���&E�1T���~t6o����űz7��=����`j�TI�4���4���dĬ:	�N��Y�^3�ׯ�ޕ�Gi�*^�j/>�+і��� KXP�x�u���A7�έ�/�m�;/svSĂ�`��Gca
%9��ƣC{cw?֮܏��_\^����bL?},z+�8��*B;�����񔠗���^_�ҵ&�5L�5�F��J�ߕ\)}����8����ƧzΎ!v!z����`l��#��V4�������BU z��5�TZ�����F=�(@G��(�	�����!�L�ͩXU^�Z
�*E�	֠��VB�]2Ӑ�K��������9�bW��f@K���i��y���h���<)��m�;���Q������ �o]�<�#�5�z��;�N����<Rٴ��\� PDJwj8� 3�"��)�^ĳ?���y��EA��[�7�#׺��Ν�՘����13�#=Z��PZ#ʱ`�d����=xh�gs�}��t)S6I��*mi-��Q�xU�X��Bv���O9'����,>u���2�\���:�$S���Q�iHSh���'�����K�8]�Q�F��ϵzUE�j�as���m�Ѻ(^G�����aԏO�`�tc���64�\vQ0�)���=d�T�KQ���N�t������j�b����J�i�Z�G�z�˨݇qvp����,�I+�(=��=���b���
��JE���
�CX��zG����/����1�}}3^��}��GЂ��]���a|��Z�ʰ4ĝI]6�P셐p�却	 �D���@Cv���5��?Ww�qK`w�0v�}�%�m<���=�m�pV�C��9ш����~36�]նk[;qcm=���q�{/\�o>;���V�s��Y �۩;$��mwe6��2�V@ڢ��L\�圄���s+z�7bnz:�<U<�r���L`-����s(h����fO��.#�~<w�@��@r����Lc~:��0%ڜ�s�i�J�ZX��"�jm)�Z�7��$,���0���F<�"����-���p3 S��5��`�B����č�v��<��{X\o��ۅ�a;{�e��zKɝ.h@Z�=
���7BI9>j�)7�Is��t�l���`x����=�?	Z��Q0xly��q%ù ĕ}�(�*iܜ���z�����UZt_}��e �0b�Qnj9 ݀�P+��Y�T�["\�I��7�q[�A�Za���g#�I��s���KQ�x�
Iv�3�N��g�,g��(R�B�
0�>�������-�:<2B��p@Zīo��k�+(	.�P�MUI;�e��-�Q��+�ȠҚ�ҵ��X�t� �QD�4�vF���VA�+� 	�^GN�|Qa�5�Z�I�	Ov���Z��6���AU��x\�$]L�,w��G/��,=�%���A�ƓF�2���
��ci� x�`eq�#y���1}S�;�&M�.a:���.�Ԑ��:D�0e�Ņ�����4 `J g]dCs�퉸�;�{��ޞ�	�c�/�f�k���ש��j���M�Q0���Wc�=;�r�p��lPF-��Tb}��-��.�܅�J� �p�E�(-�b���DM����\T%�m�� �I������!�GN�d	�K"�L"�yA^�Q�K7�硛�p�#<����7���h���A%~�B#~�#Oōý�O��bܿ��o��b��J���[����'�t��
{��q'�^r�����Mt�"B��j9ܟouvO��hc'(������h ��xE�r4۝X�݋5���Al�c�vo�w��s�m@h��H�k�� ��f@����4�tT�>�]
�z�ZG* �lS�}�w_���^���X|䙘=y)�tֈ�j��V�F!�qͼÐx�N3�g�&��aD��'���u�UvN��1o����p�~�&&0�r���i[�|1 ���J�*���Mp� qo0=
���<���a�\
a���?��4��6�b��{1�X�� ���p��4���?;G{T�:��u�Xx}�:Z	����cC`v)�~ֆQEq��x�>��)�Ji"��v�E�׊��œN��6\� vSx��B	� (��]�_����.7P +�1���((�0^{�=<���z��z���g ��ʦ���(�\=s(<R�,D1
%�>�a�����4�!���M���2s�I^�r�kr�d��B�R7?^�#e�m�刂O���.�}�����3�)�@�b��nI�Qr;&���ym����;-���i�c3љ�a�T0�O/jk/Jx����n�W�<��	��l����Ώ�ӎ�q����G�\$����u��!^I�{�]>7�8{c^{�~�ϋg���~H(:��>��39i]mYx�YL�ϔYy�;�*>5�T��g��\�EۊU���K㤡�3`�Y�H����#dV�"�9�I�^�Q���ڌ#��\��Zx0�C�Ѩ)d�C�v9��n���\�K���"-�j\��-��R/G ���sn�N�n���$�uɒ�G�R�����C��{>��D�a�}�W�!��$r(���Y.79�S����>{8ۃяn������;߸��V*�s��>���v���W~��b	S~b�E T�M��� �|��g"�M7nshA��u_@�X�C�T"ڞN�z��d��~�L�b�ހ�E�Lǀ���xLxj[�(!���]����-t�P��� `�A.g�Eŉ�z��f�vPf�B���ac�j��$00�!�88�݈Z�]��Ec~!:�~-,�ݽn��&_c��(V�:�.-�T
7�N�>�C�S��$�k��T�n��N��F��Ѿ.=�l~ó��!9�6w�����w!�;UT ,�½������fͱd����?p!Pz���N���E_���i,�:�R	>ub9���*�6a�Ufx��Π�)�d���j���"K�ⱄ+x�A��xD�0�վ"2��e��])���Oz~���qowB��#2/�&�pj��`�қ�F��C�aC��	��Q�f�1�Ed�'JK�
=,`������ѹM��HH�<�{)�h�
�Ib@Iڥ�����{C
�ߡ����Q���e���X��N��	��ޓ�P(>��*2��CaD~�B��ęe@*��P!�5��v�X���jT�aϡ�����h~��D�l���N~��=�n~�RFa5b��q���w.<@�d�XvR�N���q{�%� ��� S��m5ϑ��s]>�<����VH_���,Ī2�)�����)��+�Đ�'���)L��ϋ�'��.senAQ��^�9���T.*G�Q@m�8������g� 䨂�&p�o�D�^"2R�Q#B)`�v��|j-<=L�>=dw�	�W��sEN4�2�h�W��]��T�����6n��N�B{0��q�@�(�3�t&�\�W�Cy6F�O;��nnǛx@}_&�R|l~*�p<�{����{����X��!ֳ#,�x�E�@<�,�}�@~�Z):[=e��(.a	�t'� &q/'����s��֝a\�ދ7�w�u׺���^ܹ1����f���i���P�۩���<ϰ��h�����]]���l�����=���Z!Z�z®R*V��B`�`��ꍨ�,�
��/b!k�+���b�?����vz$%����l��%���.���♸��I���i޻�5��Il޴��d��A���\���;�KܦU�6�[iK1�F��vr
o�D��Y,�	�lOh�:W  ��IDAT�p����8S��J,b��po]�0L��	Q�l�A/�J:Gfr8�z����)x��KO<!��C��]�l��&�����$�I����ԭ7Y&� @��T�'���|q��g�ގ�S�^��$��B*U��գ(�4xN�)����,�R
!��1V/��%�&e�E�t\I�B�h�ߑ2V��СLdzb��$��փ?j;M���9酳@:�>£}��B�k�e����sڑ[H�'�E��$��+�5Kj} 3�B�i���5-�L�����H1�!�.pe_ʃ)gIA�ζp!9I�&y'�x�a:���N��a�č핾��8[f�*��9�Ƈ7c�ä*���tVF�_&��ɦ�u��R\N�&œs�u;�ݠ��MM	%b�s���$��O��F"�2����|#&�c���Y��	��f9c|���w����=lmw��T<6�X�i\0����9�6N3�L���T/�1?����_���~7���L*\�������kw� �]S�!�+�E9�* ��������S ����2�y���:؀q��1jW�96ߡi� }@Ym΄QDu���YR���)�2�+6�֭����L/̣8t6��Z���GL�V��B�+��Q���C�� ��`��/k�ҧ�}�s%ͱ���
+<�n�ы�ʇk�STG�Q�i�	W���ٸl��?-`ې�]�y��
OlN���ga��kR����
�:�1M]��8җ�>�����Q�8���a� 8��wi�N�π�9p������I/h�)\�ķ�NV��DͿ���o�����X��X���(H�s���2��v��bl�*L�26��܏��uY 83i����a�p��E�dr'��|�$~�?ӓ\C�k?O��D
v����u�v�C*n�㵟.��!�U�t��:��}��*�2�����5Bk"�S���)���L�`rk$�r��R�K?*)q��m|QP�\�9�@s��Q�"�z��q��o�{�0�21�S,#�]�?�+��¸���;�ht~�H�	}P�k�\���68�sx#��n���q�^(��p,s\��~<�Q�6��G�a����;�(�Ҏ���3�pqD{�֣��S�|J��Q��*�\:�yB�A�2�͜A���s5�:dd��D���n{�/��lb��y�b�_�Q�����Cw�m	��y��n���^ZI�s������w����x�N]�+�H4��L�Y/9��L�vo�����_y3~�k�5c�P�?wq&~��;{�|�������0�)�wlꩆ�P��A�\d+�E��D�6]��D������g�L\��
��A� �*���,�ͭ�غ{�jC
MV���!i9K���a��}1��d^��ɼtZ����JN�d>BZҖ�0su��7�O�%|'�i'�k�"x���F�a0S��, :�1j���I`#����UP�N�bZ~��~�cl94��p	���)�߼�e]]U��r������:�	���B#4R9Q��R,K�E9מB5ءͤgk>���{�1\ߌ��ݨ���4S���C�+KQ]ZW�{L<4Q�yח�:�!������VP)q��W(`W��Hx�+h��v��L���^�~�#9LC&�þ*�";x�,.Ef�z��ף�T��L9��G�?}W5;1�@t.]���(�3E0Q�e �?���4� 	�и���?��x�m�q9=�׾G�3g��u�H��gY�FH��~����^���&,"�ɏ���Æۭ�ﶣ���s�*���g�R�

��Q� _��Y��t�M8I�<M�vn���^3����t1�-W�v|�{.��FtKU�dw��.ꘔ���[m�p*��]qb�L�q*���C���#�7�����Wp�F	"�yp��=r���$Y�V��b=y�&
X�Ϟ���R��Uw6���)�f�5K�:*������\�;��O��p7k\�]y�aR`v�&�ZN��gx_X�J�kN���/qmD惢-I���sb�	�|㍢�U�:L�Z�M������3C*�B���f�t��h�P>����+W���-Nş�8�cOƝ���;�z)��C�(�i,�*��/RV#���/�I�
R	�F	3i�S��b0��m�H� �q�eߪ^���k.���M�*!�U��E��^�X�ZZx�}���H����V�Đ��J�8'mJA��'����
��N�q�~L�Rw���䰛>�ˤ�Fe˯BV�£?�B�C}"q~W�!@]������ ��E8���UQ*��1� �KK�V�;���ISXξ���t�6;�o]���
�eg_J( g�
���A��6b
E䇱|I��$(� T>���9��T�҅#�ѿ�^�M��7��~Ch�|�QN.:P��#�7�ݒ����z�)(�_5�N�bTA{
z�O�i�FY��H��ڬ�A+K�����S�@���A$Q^Z�
!`P!:�'��4�3x� ��%��&2'��Ԣ-�s�|(6�+_��P�����yA`)���)��j�m�Q�g��P/8z��;����jGg���&^�[G�A^&��uPU��S�.P��Lt���m����[G��܎ҝ=��!I�j��sF�./E�1�V׹/ڒ�lL�	3'�/�P�����m*�E{=�š�����<7��/]���Q��G�֭�/x߃���X��3�v|�"�7����K<�N�d���:M�L�_
:����k�g$�7	@1�g�����k�ǁ�S.eޜ������'�x��y��_�������U���Sbq·���N
�C"��G��  ��袡�x=(��/r����v��?�����j\<�ۇ�����o�p���hHUA!r�:������~�a�mF�+��UXU\�z�R�\���y�8v!�N�d����
��c��2^Mef�v`���i�����P;�@�K�$I��=>�`�TA��u^�K�BH��NQ�q��B��m��(�\���7�(!��
9������hI��<g��OB,�8y?�D����r���twE&is\��",mᖼ��u��so��{k�Tz@�{(�i�fy�H�`�<F�u(���?r�
/���]��l��btU��������e��*�b�9��%��'�<��0Ma�d*�:J�6����ʵ��тO�y��x����:N`H�K���}��'��9��	R���D\RU�V2k��y��&\*���4����G$�1�Q~�����d�>R�poH �>Q�G�&+������a�}A�Opֻt�����͕�v�Ar�>�_�ęBS�?���S�zrVq�b�r����v)��L�Xf��I���Q�r"'1�"i�QK8W�]��ϸ��G��"��)����xa7��O� �|��g\X�8���ѝ���(-�Az���2�e�q���'i�%}����".�!���Y�i���I3^KO�8z!N�G�0���r���t�C� "� N�ˡ�	gQ����]�{�#E����i˴<n,�����%�� ri>�pC���e���B�a�1��/|��:��k(��n,��iL�c�x��rlS�woމ��Ӫuyg!D���|+�ȹ4�4D�R2�9���{���x�5Zs�_	/�OpXfO�R��Z%S-�ʵI��y�I'A3�ڱe'���U��$h �IR�hzZ	�)\�N��O�'���`=�c%���EM�k�P?����3�����d���T\\-�{�؄�|m$')�B��˟[��k�9	�^_�ErR�Sq&�L�hĚ���$\�=𨆩&���_�s�w�(7���Z�b(�D�˖�;ƄH)��P����ʗ/!�}��`��'����7`��iE�{Hq�Ź�>@���*�2Uo��"^ʠ���o��=�r2�k�V�g|.w�ق"��e�4�JR��4�����E1BP*��`CW�"	�<j;׍��A�}W7�{ܓ��c�{? ~@9�B�z�br�x���+��<k�i��~�;nn9e=���O~a���kv(xL�f޼nu�:g:7
��y�
�p���k �I_�W�d_�7�� ���1W�.�F:�J��*��.�(�3��r�6�9�@>w(HC��9��l�,mdGQ���5=诀��y]Z�'�I��H���NX���"C���(g��k��MXԟ��2��G^'�2�?�2�0�
�Q,�l|$,���c����u��g�P��`r&?
�'GÚ�|��W�QоG	;"c��C* ��r�))�h�m*�R�[m�M܌�7�j4�K�|r�GIc!>W�8?&NKJ�O������_\�k�7�n�z>2]m"_�Ņ������w�߇
fϹ
�O(,�YTb:� ��_��H�P�M�e����N�磌��2�}4��R)h�r8��%f�/|fq�UbG�ڲ����;�ZiZ	Z�U�b�>��d���1�V�sJ��{��m�n3Q)�	���������������šh��WչzN8/䋦������	Et�B��q��B��²(Z�!��:nd������V1�ΈDm���Q!��Az<�4i����u�B��3I8I�0Ǩ���V�o��x����'�4
l�G~f���t�!�R������p]������+���vQ)'�����P&ڤە��<[�L`�}�3� ���^��~���w��V��}�?�����#�{�>+��{( ��1�g���k�vt��3n�K0�~+�0+�3?����&�ee�xV�-졐�Q@�%ݭVtI�q�M�����}�8�,��E^�Ab*zw�w�#H�
M��9�	��t�B$;��<�ݎ��T@�tU������L�gzǹҲ}� �]�1�!=�p��$�<���C|�]
�▤�
�ʕ2�2�N���;E�"�'��f����6{?�{pU�'�O�����ϼ�~\�I����Iwc��CZ*�y>h�ܢY�����N#1�-~	lV./��F��� 
	�gv�g��d>�#hsh��,���{C�'Q�ɲ
R�p],8@^/�_�,8�a�$"��ό;|�k�ׯ�Ǜz>Μ#T[(ǉչ�m���z�D(scw��zd�C<Yl^s�!l�\K����)������\<�R��	���GA��=�yA�]����Mal�*.��c�}:�a.�ȳK耾�:�ֱA����s�=�׭{/\�X�N�N�q{��C�:q��������R�VZS�X.w��R\��sF�������Ș~�A�#���:�0�)�U��k���}p?�w0'D��_*�v�s�\��^�O������s�a3f��Q�i����ɋ�:�dJ��J�3���g
�;�Lg�a�\��U.��̭�q�M�գd��Ez9�FOT�����|�x�6p�*��������r(�G��s�rTZa"��|���W$��y�	�;�'⁐��9n����lG�~v�������_�k���E[���j�mH�� LZ�?��4�W�������@<)�>��x�� �܃�0�:�A�'�����Ír�~��(7i�]�0G�����,�����s�k���XjLũ�阞�R�(:Ѕ}�CN����6P�(7R��	���S\�R6���t��ԥ7���9�j��2Jʕ{z�}d�;����� �y�wGO�0eѷ�L(<ARN�Ȑ��?�I��g6ռ)����q^e���x�W"g��H[�J���q��H\� ǹTy�J�;Q6�W�K1LJK���W�m�d�9^�0\ѕ|m}
L����l���=��eZ�\���y�b|��PomKڐ��^qd`�|�H��:Y�娈��2*�vK��_��}���]]��Ww���M�c�q��jt�Ŀs�n9�Z��2g�T��Ķ�IR�`��4<�
R`�����9!�F��P~�s�[v U@-��Bk�=��&^�vH�S��Õo����M={�&�X��"�G�tQ"<���{:z
�"v��&���A�{���}���c��i����B�w��5�;�rݳ>w8܋E�@���}�޺�׶��K�|��wm��
L��:��ď�A"�}x{�߈�7���0}-�Ӌ���!:p�����
�	|��8ܸ�e��3�XZ^�)?1Q��	Y�0
������;��3�B��L'��u�nt�ߋ���T����pQP$�mR�X�C@O��g����BdZ��������uA?9�2VP��vJ4'��G�K]
y�^�HDb�,UR�8�~��EY�We�C��F�4,��٩/�KN��Gz��V��{.n��ط�R$�-z���їz��,�o2��^埸�`2�FXmC��W@[v�y$�������	lqA=���);���⊼���??�x�����Z%v�;��}��9�̠� |ר��҈3�va��zݹ�y3۪��s�
X�գ_��u�7���K���.���
��$�ܣ��}H��yM�}}�qb҃%%>��ś0���ه��(yp6�2��Y��(��l�q_@����8)$eV�y�etw�)��,tH���H���BfUd�Gzy�����G�:��,*k�kq�Qdd���QZ���K��y��d[�g;�$�m��w�ݬ�4�I��S3]!xƜ	dF���b���/��m�W�n��k;T(b{t�O�� vo���<�@���eM��1��'c�I���.I��T��u|[�õo�;��d=��
I��D��'��s�H�������k���n��1�m�-�Fw?ۭ~z��� ݏ����so�h�p��k{����؏�z3:��ѿG�u�٢�M�wH�����Xu� �P����;q��w�l�囻q��~�!�V����u�ߕfP�䀶`�%q�n����%ؼw%��;J����?���Q�ΑV!oo��������X���G7��&f��(f���.vv�A�@�y-��c���¥�@n�c��غ�hݽ����Z�j��A;���c�Urx��a�0��f��$_"&��ι2U�t�Ⱥ���s59}�ۡ��&/rHG���KI���Vru�8���2����b�RH� 3.�N!O�H��W�[(�#!�٠²."=(�xB��%�s���|x���a��0�.K�n�i0�?�ѵ*�:sd��L�E�\c�8�Ó�CwU���&ca����j��d�l����tJ�iqcA������U0�����LMe�|ޏ/��3=K�T���S}u�����`Xf��ۛm1�F� ��6^�֣h#�$n�1��W��:m���@{�=B��aYe��p]�i-��č�=�)�N���D���p\|ﷂ®��(���~*�d9
kB��X��D,K
� �Ko�G�
�g949�\`&ʣh�m?�E�r�K^P!��<o&"$m[�N��$<\ȼ��!��&�L�r?�2�4���˿���k(�+�w>PL��B-N���A����Bƹs*��j�<�# �; ,�N���I"P�������Cz8m[�C���0~j�/�f��]Q��WGA��vZOx"(�@��%�A �cc/J�K[m·�׵�*����u��X��<���כ o���'%|��h�<*�ݬg�bm���XkZ��z���ڍ7��v�̱w���eo��Й�h�+ +���
���^k?���d���q70=��8�c�"(�EHa@~YԾp��	����tz�]��2�ޏ����1[@RH�~�ˇ��bk�J�Ř�nGcf)jK+Qr�b,Z߇�X=rl�V7'N[0P�A�J�Q�_Ct�Iik9w+��l�Pd92��L>o����$�J�^'��8�U���8@� ��ud����o�Ց�z�V�Fi��5�u��2���HiT�������F�"O�Z��0�ϭ?=_aI�dOd[�.�P�i,�Ao��+/��	%�Fq���\Y��xJ9�1���W�ok��C�҈s�8-Z�6Z�u�����
|�w��r�S��ǹ�%�)Q�@��|n�D��&9SUT��l=�x_m��v)pB=�d>���E(��b9��G1zO��(dGJ �@�Gىk�>�ȴ��u�?Q'!�㼔��G�QĊ'i(���ȫT�G�։��a,L���p'f*-���&eW9F��[���cvu� "s�%AO'�o�9�

x�o�N�
Tx���g���E<�4>#��S������E�8��^�C&�(i�r��?�}"$�|�T>x>{�x>�q�ރ�nx>������t4��x�a�z�T%��lkP����R�~���s)0�і��殲��wD���iU����Xwӹ@�`w�ˉ)W���w����ߍѝ5��N�_pt,=Wu������ެ<����@S���^I���`0�C� 8�1���9!>@p� En���\af�I}%����x��]�&
�t+�Q���K��68)�p;,�@}%w��X�Z�DL�s�X���wi�7�e|n�v�PLK:����T��.k��'QN�c���$��mqr��"��?��o��mҝ,����'���V���^�#��P�ݻ9T@�T��ĨÏ���ԒYZАLUv�	�fgߐt�C^q�n��	���yRAI	s���3���*.�E%א��}) �i�G/��>E���QW�b.�-���a$��r��ϼO��0�U�����ʳ��L��Y��#c��*ز���Y�G��W��N`~C&�� �Y�@<��?�܃�˓�^�� }��B�\�G_��P�l��_���a9���m��ݹ{ �[J�|�P|�]Q�15?sQ��|��B�x �-ɶy�8��PqU\q �4m�R� OdK匊'=N�2��i�X`Q~��(J(N����菣���0s�0x�R�sD�N�z���9Vڊ������Z��wby[�W��G"eƂ6������M�q*�lN68�9�/q7���By�g�g��d|��#�0~^�9n�7*�s���t�v���
�^W��	��#gF�:��hn6&���Q>o���5�h�|���q�(�����@��c�gd`W��d
D��>;d�u?c�[� u��s�^N) B�%��QV��w�_�t��F�f��Rk�F�"��gsgA���}�k���Ɇ�"L�E�%B�7ؕ��0J3���]a8'>�0���`f�(��x�
�)�u%�}����Y~v-u��9[`O�\�F��3x%\'��L�
0_��r	j��镘Y>����_�!M2�M�Tr�mUAәS���`mbM�O.�ւ-W`/�Kb��g2��2�?�J#�:h{��gkK(�SQ�;I;��H@�*-��+u�\=��)��49��PH
�έhj �\Y��;E�Kɍ����P�Ͽ�����&�/1H|��m��VL'�]^��o��ނ8�����!{��@�(��L�qن�?�C�MK�4Y�m����6����'�S`�L�_�vSR�If~��ih�^쑠4�XH�Cq�9� ՝my��zip������\6����40ra�!!�M�S��\É�Qc�Ha���C�0}hCcԍf]姑��i����11;����pQ�!��R�E���~C���+Օ�H5N4:�Tb��m�x�̴�WƊX�+p$m��y_\x�0����&ɽ#�9��nó���b�ލs�X:x;^�~l��R��6��L=�_���wO��\�Gy�(9��Ǯm�,G�E$��h+�(�Ǝ3PG����w>�D������G�v��� ���3����4*l��P���+d��l�[��������k�߸�P�?~6>���h��������a���`u���qG�z��p ⷰ�� �b 5� @�7@��J�҈'����L�f0` �}WB9���]�s{;�~��h�t<9�ZW���C�qb!8�DYGouG]c���qj�й�����Ĕ{��$?xU�	�]�>-a���n\���V
���(��dr���C���qok+n�ߏVEz,N]8�.��Kx�0�+��M�rG�� �)�b�}L� p�t��rɉKACx�'	~Y�X�K�%,Zw�	I�T�V���i_�4l�T�&�筃�+c��^[ǯ�h����UA��;P�#��Lg}3bc+��_�t�*\�bϪ���,,� O�/�:\�vߵAͦ ;h�����n3&���C�ؗ�p�JE���T�ˁ�/D�!OE�>�kg����2��<�{�d#��D��g����?��`6��������<�b^�(,z�%��m���N�,CSd�S!�ɲ��yQ�y�ĸ5����]�Rs��$ʀ���1FX}��U��;m�H?2ځ����y��.eP��X�!�4J��
�km�3'�"N,�&
m_��<����Q��hf�D5�/���q�7���Sf �$ě��/���q�p"�x��rH���%RIԑ���ľ��卣��v�83����BS_~�E ������x���ZזT�mz���o-9�6(�:݉K�x��S׾���7�Ƶ�8=���|0���x�U�?ؙ���j[�b�C�H�B���{@��֚ƚM#�p!]*ãHw�z���,�y��d�����{S����.n��'��;tu��4�)���Q�:��a��Ũ�
^υ�*����[�o����|Zx�g�3�>�u؋������ �8j4x
�b2�x!�Q�F��nstKF*����m��P0�I�b-8ӈ��D�=V�w]Z��_<��NǬ�����9e��{{�����[��7b��:�����;?�g�z��S?�r�am���	U�;��7A��N?~,VW��q���CkӗK&R��x�$���.#|��|�R��l��p7Ir~khc{+^�z7����7�b�5K����'�!����Ӥ
����*���Yp�,͞TLM��k�c��gZ�� ¨R8���| �B��Pԣ������t��ÉIb4hPe�̀��"�\�|��t�ȡ<�r3X��qh��O ;{�C����r�0��%5�P���1���}-���i����>��!}�nb`�|�W��{��*�G�Mp�!?.ؓXl]�Z��dSms
�"���A�_*�˿3m���eF�Dp�`j�"]�����d�Žװ��3�2-h�w��d2��'�2�R`��G&���?����4䐈<����rx�/�5�Ǝ4�;H��V�
g�a6\��.F�ӯ�6���/�A5;1�"�
������7;�Y�Ʊs�Q9�w e��q!�(�{Q����Ub��J�N���T�w�a�T>Z�6���O�rX�C|�aZn�E���� ��K�(MI�i�6���a"j�D�oQ���{|����'����r�����$��K�m�E����^��<�N<�Ќ�G�Qz�{��?�Fܼ��C���ԇ�̇?oN���l���=<��?�}ҩAz���2k)X�d<���"_�(
zLyWHr��g�2>�ִ�"˸�䣌�m�Ȥ���Z�uW�r����4����'X�_!.�|.�|ڇ������Wވ/�Vt�q��
��O��/(�߾�Bt�1Cc���Ձv�k#@z���=����>�W��&6���w5�_��'�:KKq�^�G�j�􉙸�Ԉ9�&_���F'��(�~������ߎo��c��ܥ�?���O}���v($���N$7b.�>88H!~���X��v��a���꽀+=�0;I�%1����jD�r���ڧ>�����T�A��v�n|폟����o�k�u�B|�}OG���[��J$���nQ�`h�g�c�1�} '���te�O��(��[Ӻ��P0� ��T>��?�Jf���@�Xb.�~����f�^M��+��S9?��@�c���� �+����v�ֶ����f�nPY�ӵ(�.�B��R�AG9IE�r�7��,����y� "?I�����������g'B]`*�ym{�)2f�
A!3�ش�4��NV!>-K�����Ǖt!����Z����=L8>0k.�6��Y�~�+ķI���&�p��&�AK��FH�����N)�1��[{qxK���V(�x�a�F�uhm����g��ptՂ�Q@]������w�X�W�X�u�K�>^B��yh5��M�~�O�3|�P>���g��R*��Qs*y���$J�,K�?�+p�2����KoR��������Qjm�p�m��ͨ͞���#ѫ,Ge�9�
�t��d�$"��qt���~�]�	q�=Y3�,��d_��l7.����S�����o~)n�z;N����cᙏ�먢n7b}��6�H-F#ą8w�Q�vt����7�yP!0�CdӬp%��eq����ȣ��H�?�H��8ۘ�77+�Rv�=�a�0�;;x�6(n?r��#-
��슙�<��ep��n'c�����ϵ�v�R�zyj�N,��8߻y7:�~� >K
-a�}�Fܺ��y)&�%,��X-M�,k��3O����Z�?�����}�R|��c���̩�8�R���,Y`���n^+�����-��N'��x�r�8w"fg��9(?�P.Wr�ֵ_C�����ՕXXZ�Z�0��Z��
br�;�;<�>k)�-P��t���!AtPjM�/	��AEMM\���wbw�^t��8؟�w?|<��˱�{K*�zd5�Qi��b�R���E
AbS��<�/�W� �X\��T�Q�ˑ��i����Z���OzS�/�a����3P	��&!.��Tj�i��o �}� �+���ؠӍ2�h��Z?�m��j%	�w��N%��u<�O4PX3�*}X�r�]�}WMv�����?7�1�X�/8Z/�� �r�}��L�p_lŔH�i���Bl�π	dfZ��i����8���3�r�Y�x�P���.h�X�8.� �X�ϊp_�m�yM���8��AO�2������o��d�Ɔx����������sl��Ck��H��]���V����v6c[NҰ�u����i�͙أܽ�s���J�]<'*���`�/��D��Q�pHc��t���A��LGk��"H=ߎX"P/���Z��^�r�vL㥗�1���gR���M��A�,!�)��W���z�Y����[�K�E>�L�e���;��Yk���أ'�v��خ��{��{X�ng
`�&*.ZC��j,�P�G0p��y&�#���l���zpX���x��>�/�ʂ�(�1�{]�K�QXf�p��"���L>L�����ن;|!7�����rm;���yh�'Vx6�x��zt���p ���o�U�X�T\�u�;?�Q���&����f;���X�_�܅��?�p��s���V���F� /\S�|}�W���Qt~AX�!?��.��Deה�y+��.��B�u� ��m'�WG�4����!�A`TL�QKxt����F��l���Z�����Fܹw;n߽7�܉�o����۱�܏�o��ٽb���Պ6���A\�~`Fn����x��U�m1�ۥ�ϱ��hov,C%#���%�
	��(�Mc]��&��@��{�\��H�}�C�ZD�K>��$���s�Eҙ�������5��ȧ�1	�Z�M"QBIc�*ƞ��p�B_��d~/4��_rQ��C�)�WY�h�[�m�o�c�ObPF�2ZТ[*0��J'=e��O�D�'ذ�뽍- �y#�@��,�:*�dX\)�b��>2_zM�</�>��~�lY�����U<�s��C;LV�����b��x�3p侈���uO!P�G!��#�>�Z�p���+��
���i8؇�_e��W����Q~���nl�g��c0�/��(�}��)]��ь	]_��;ϴ��:;S,8P� M�^p���)�Hq���{�HZ�:�4�ɭ�2p��3��8��!�����T0�U�_(�)6�������J��w$H<�g��%-�R��w�+'���41��cgcb�؟>w��q�[��6�R��NY�_�W0�ՍOYO�Y�!�Є�oR�� a���Ē����r�9��ʲ)ڼ���̟I�`�+j�0W���ȧ��u�>��'�j�9�_��_���~'�~��|�s��1���|Vp��g����\�6M۴j����B�ZP�VL�����@�}�b�~,>��Gⳟx4~�c�Ͽ�\|��B���نo4� ��([ek9��w�];/;�Õ:u���(#X���N+�xy-�^��}/��0GΑ�����m���"�,k+*�Z�n߽�_~#޾z=��Y�N��2��n;���c}k7��ߌ�[[q�����ո���M�>
��*e���v\�v=�o���d�X��#xh�����Fq�.�q�!�jg����<��h�K�ء>s�#_�s�h
�9[K>?Gq|i6HtE�$�f=���w�P�T���۰�U���	T�.(@ṗ��A�zn
a�۝e%�چ#�-�/���$ɝ&u�avW<�\��%�
����L]Z�|?[��e>7�użJ'��Q�ض�_��T>R��$��$_dZ�%�'H��;ƭy�T� o��T�	��٨q���� ���Nڬ��E^��TZ�d0��7�+`Y>׆�L�&��,�gG����'��Z��ޝ�d̉v[|UX/������r���,4�a`�hd�|6=-���Ŗ�P0��w�9Li;u����ӱ�����0<��͈�è��1�.������b\P�:ώȟ�f��+^'�
\rgEt�+g3� >��;?ʎ�Z=&�OD�|<�%�h� ��&�N��sTW���,�E��1�I��4�f����<Lm,�}��dky>�+K�9��-�~�:i5"�����(-��sH�,�4B!����0	nQ�=�� ����6�2����,�?��#��M.��ޗ��hW�K^r8e� ��48"[?��/��T>_��Y(�C�X��/��91�c�/��:�$�v�M�e�(� ��GH�rK-*�Oć���+�6���O�s�S�riT��5��1��h��B��HUG.�F�8�QQ�������v/�{���8�TG W �a����4�{qx���X�C���W㏿����˯���Ǣ�*���X���q���F��kw�������s��뛝��c+q���XZX�R�[D�q��7�ֽ��~8���R��p<��q0�0-�Kh��N����*:�{eQz6>�g4 �y�U!��C5��$M<5'�(�
z�<\� Ѩ�<��8_����Pd^w�]�x�#�" #��ז���1�1���I!o�6)����h�Um�N�I�_M�Y�"�Ҥ˶������}�;��+%
ծ'����i�e����J&q3Ns�Rf1LA���X��1Tx�ܓ�t�7�1��0������c�C�SL��ض���r��])���6�RF�xun#˵<�e�������⧡�����Y��#���)ǽC:k�,NT�(n�C�P�8>#��If�N]1���ܭ�>��"@\1��;�x�'yN�y�|�(�Q��i��3���C4��+d�h��T(�O�6σ2����)���@/��޶$�w��1�Z�#�ڣj�*Ǣ=����$�8*f�N�C�d��/DT(QC]֓�q)��1EҔa��_z���� ^�7��
���_%�tz5<z����b�%.��}�i�Ges��yO�����CX,����� ��o|]\ej�&^����W6i8��tح��'�Mp��P<	XR`iM��g&&��+����f/�~m3�vshı����qry:W}��z�� kȽ&@�j7LlQ�/��������G���/�/>��G�̱���),��_zh�<@�Ey����AIO)ILR��?�]��fFq��t<sj1�85�¤N���;� �<h���Flnm���z\�r9��x+6����7���~|��/�u����ә�阡=~k�Q��K�3(�ju��0��VTa���h,��C���c'O���4J�w:������cc���|��Z���lla��+smMz�_�9� �<۩���(�B����w9��[���3�C-�8F���M��.��N����P| �ٌ�A����&���m�;(쮁��>�{��v�����>xp2R/K����Lx�T������� @쿧=*��@T/�D�U^�.XQ�-!�]έR=�la
*,���ܧ՜U�Cw�H�$�s
~��^��N%{`�i��.ھT�K�-�xw�&��s��>ew�<Iظ���t��y���{���?~�䬻��{]��H[+��^��[.�O�����bL9w�^zy���2߁��3�Ct�b+8V���y ⻔���fг�a%hw*��L��L=�u�7�����5FG-�hi�"\y�G���O��K�]�|���}���Z#M}f**�uxb���Nw%�� 9{���n�0yd��(N��#��|lY����ৣ3xZ�|mp8�P�L�&�{><Ge�����<R�x?�K��!�%��4()��P�x7CW�h{���ٗ���Hk����N�x,��"��? !+6o�\����
�({&�91f�,�8��e�$���u��+yڵe��GA`�eĥ�'��������xw7��/��菮F{B����_���;�;<�'�}#:��	�@ٌv�h�B$~���r<wv).]��?��S���^����V�8ޙ�j�5J�`�����tE�s咟@nSv�ꆦ
�\n��FZmS�BX�7i4�w�^����dNvZv&�����N�mm�>Z�����w�Q�^A/n���l�RWO�gO��#����/ł�U��&�P ubo� �w��QAA-�.���'��3�X"ZY��������?���_�T}2&��O}ꉘ;*�&k�&8Hf�N���
Fe��Y��������ѩ2���"+7��˾-�Ksm-�(�
��Lz���[�:�:������8��(�R)�}֧�1���'��� �R��O�16�@��up���(�m�4�2��@���7�(��J����L@��S����2G��z~�u�:�U.~ �g�����T�Fh�r�Bq��F�:T�8?���\�簤C�WYKU��T��w�^�.���}bG�0A���֣����>���#��A(��E(��#i�d�:�<��|L�U�'��Q�M�v����?@9�݈��NL����Q���[���رr����X���j5�hɡ��m�Co���>�	oi8�U�2���K+Ѹ�7P$7���<��Sw��ͯL�ܹ�w�^@G�#��AA y)t� J>).3��6%�E4�'�J&
���v�ˮM��h0�x�Ka��(��h��#V�Eo��$o�ݾ)�O�S\�!���)��LV(E�#$�Q��л�M�\(���efJ�D�-&۞Wҍ�V,	,��%�h�r�����<�ЀȢ�'��,�T����o�-�D>+^Ƥi� o֭��ϣ~�[����&-B�|�'�i�_�TҸ<�C@&��\���S�w��ڌ/����_;:�ť�j��ř�ȓ'�m����Rt�B<�t��ڥ�=��fc⑹���]��ӏ���c��s:���'�)持Ih8�8����a�7�w����`�a�����	F�B<ZE2�+�V�cya:W�C.
9�D׼�N�]��god��51yv��x?7���{Y�ʭ�e)�+x}g��G�'���梁%�'�p�;(�C�[]<++�q��1����i��qM������_�� ���Oǹ�>+��~e���oB��!���I�N��M�?�(`�v�'�0�1䛣����v1Ds���kQ�ވ��]�S�I3���� |���!�����<5t�����
��*15�О)�;��V���,�\����0� �drTI�2�H�|����:���@vc�V�X�Ԑ�(ȴ�T:9G�?)��
���$�p�x;DȊ�$��F�s�"���B��'��k�Ɉ��}/,���L|��T�\��qje>�0�޼�M,y���[�k��a�B�P�����j8� x9.�@�n\1�����	�֯푞���by*���	�()��� .���c@,��f�Q_����|�f��N��v�+��@c���\&{c-b�9�S��0~*���^�/��r9�fc�4wQJ��t�{k=J��1��.��(�Ņ�8ua)�V�0�:��k��z���F��痧b�u��1�BE_N�/a�W,x�?�d����^R�仅җ�V��X�H�)y�{M9b`yI:��*G�|��EeG����_�y�||d�2�Ϡ?��w����Ln�B$l��L�4�q���xy �%&�/���$I��r������h/��[�:��\>�#�o��\�����*~�Գd���:��A�w��g�����)HEv�9���(����R���O�����x{��}e#n]�ƅ�	�S�.���+ :�x�f�uEO�x�V��c��k>������ǧ_��˵h�λ�Y��!���(���!̷��$��X�/vBQ!&�1�KYS��1@H��<L�r�4nq�C4ba���g8�s(%�7�Ѯ��0��Vj࡜ַ2jnn6f�
��ZxO����6�   ,_@�/�b�7313�u�yfa)*�i�06[-��sė�`+UB�߸_�{����ct~>s(�jZC� _��TbM�ɡ"��e��^Y���R�����X��<�|�I����Y�SAOm�ӌ���ypYs�`�䙤��N;��p�H��#�s��1���efx�ȝ*�x�
X%�mu8cMKdx4�xb��ZYC<*'�i8��K~iӡ2 O�����e^����O���Mv-�Ĥ}E_8Tg�%N���L�5�D���r'��I�'b�v+�����z͘�\��t/j�U�3�h��T+>�a��^������X���z̏cq�0fK{1;a�=���F]t�����z��]v1�|I3?G�wxz0h!�X���ZPv#�ޏ� �a%؟6j��yO����J�G4Ԯ��o����S~��R�+)����v�sҗ��h��)V���.����E}n&Z(Wl*+�*i��2�¼V+��B=&1Ui������[͘�t�֘���:�|�4�J�#�؟��8��A��9�p�%�0����H��IAN� �[���]2�'h�6k���6ϖI\k+��g�fE��>�~����xd|���+;�gy��qV��+TR�FF��*������^z.Q!�
8���p%y��P�x�06�y~����b|��:��T��5,���R����F����W����i��W���/���į]��R��&��ŉ�t|%�T��7�Fw���#��h�h<<���_��񞇗b��.AT� e66���%�w?�M�vo�>�w��n�L+�:�:fkx�--�P����k��X���c�Wczv፰A�8��� ´
2�R1!�t%燴�OO��LO�4
D���HWq<�k���5��J�ꍘ�������s�Q�������p����ǄP��c�D��ٌ����`D�N<���Q_Z�.^���ss�K�ӧ�^���^��0�Q����� ���ߏ6�w���}s?�:os�3�uT��C�ڊ�6g�8����
e?ʔW�w\�O(��軸՝�^�Z[�]v�����A?�G����:��bt��׎��&�1�<�.��
\a��x���r����S�i�;6qϵ�/��~��If��m_W����'��ۘ١&}ex�s5�j�� �9�$(��(��섹Ln��A<Tߏ��ͨt����V��v�{[1�]���6��ߢ�>ۍ���N�Z��ӫ`3�ݼ͵��>\���<��ܨ��^L׻ф�wm���$�t��/���^@����pBϡ8�%%>�+6P4nǄ%9L� ڗN�ِ��o�W!��$�}�mzG���'��,����C�a	�s%��-R�OT&
#�]�����t�gcA�Mڑ
�az��ص ���U,�(c$��F4�-~T>���7��&���r�u����Sv؏��sK�<��� �R�{m�w�j�<�ʩ�خ���!�R� g�� *���g���g{
�B:k�4ɵu{x{4���9�2Z�'t֝�ič��2�G����r�D�b�����ƙ�������SQ�o^��(���R���d���A0�GA9,[<��HW�%�a�x�G�<<K�Z7���tL�����;;���(����(�yx��:��[߾|'��F��4/��?��s������E����f��C�9c���V;�6���N��tu��0���da�A�/t��:h"����+�ϹE^ߘB��J5���h���Z'f���b��m�`�8�p��b��[�7fP� �U\���g����j��n�4^��T@33�Q���*WsABX�7�e�O�j��݌��?�O
�/]��cQ_����8����o��n�-X��:̹x��OeԊ��r&��t����lơM��8�>���DE0w�M��]�bG/
��*���������Utݭh��
�M[{t48)=t:�|����O�+�̟�`�䧟���I������s0D�:x���8�q����e؃F5Z�?�^�����UR�F��_���!��N=$�����!0߇��dD�������=�)���\D��ֺ�NOyX�S�La�3w��O��R�^t6߈�{oD��~tע���z�.p�� |5Q�(�3���ݸw�Z\}뵸{�M�[ r���6P��q�o�I������ ��
���P�$mW��Kߏ���R5�7�	@��n��� @�N��s����偰�o)q=�Q�0��+u(H+.EG����om���h�!��=�@(���J�(�u��K���w�d����ˡ�e��Uť�����K�#=-L2���O(h�ɣ~*��$�#��ӓ�P��[��|�EZЃK��T4ye���� oC�
�����棠璒��9�6V:�|��}Gi
�dY�+dYO�������2�28���	@^�s8\xtg�,�z�+��!���l[��wtXBzL��;���:j��+�卧��b1����|��w��������s����~J_��R�{i&�����R��s�V��j�_���{>��&�ϭ=�JAP��pά�s�Է_��p�@�K1zx>��'�����-�Hč� ����^륍U�S�`���\���A�����.
�"އ�v�0i�rj�.�>@�t	5����K�hW��x�z= ��S;�q\(Ux�;:�9*xCxD"���2"|ɱ�qND�Je*�k6(�94רK�2Ki��-�
��\���o�o����L\���(�|�� ���r���Cwk7?QÚ,�J�N�8�*Xک��W�����=�l��\� qQH�|z�x�e(_&m��C:} �˳���3���~������cerf~|��x�]�Fi������O}:~�?��g���c�ѧ.ŉ�'���뱉ǵy�k]O�wR��J��8�2�ݹ�=��e����6P�5گa?��F�v��XߊI��?�aYu�'�����X��]��sF�
P������Bm���Ei"2��c �e�	ʜ,�G-���[x��)�I?L�*Ŏ���
F8������ߣ�]��m�*2~5e#Ji���p�������F-&�x�9~�p��(����}�z(�B�8�8t/;���f��Gx��ѿ���-�#+���K$j�����ל�A��d������L9�g����hMV��re"N�L���� W�_��gG Յ��/@����Z�@��U��^��:ɡI� ���ZL���j&�|F4�W�i�Wۘ.�̼/�����92���Gs$B9f�)��cI�����e*	�T��gȳ�T,*bp5	=�l�̽�r7v�X��Лuw��������wYM֘���~���<J`ZOF�<�Pd�Zz�����ezQ\^`����T<suߧT�a���4X�� �fϬBj�g����G�&/�1�	�/z�y��+O��j��m>�h�)�U>x>��V��卸{� 2�YB���@8���w������w.��O<�=�Q��Z;%6��ˢ]9�m���|���qS��-�1nZko?��wc�w�%�r�<�|�`��v�%�ՕcXO�����ة�|˺��v9j*~��uI����R��u%xV+��Z�a���
����|~.����m�ɫ���M��sG.�aɗ+*�=���F5��+z4~�;ߏ/��o ����U�c��Ʃz>�-�9_R�����KI"���$=��1����V���b��&7��G�kA���P%�[����19L�Gݴ�O�U�C���=q�_���A��vQ,,��cgO�O~���g?���������+9I%����(^���� �!%���$r�\Eؽ��\��w��w�?��5,䍨t������io��D+޵҈�+0�^Z���-��s��5�j�a4]�؇�$�b5��W��z��x,�=�����INLO��S���s'⩧W��I�a� Z�w���V1�00c�6�ЯSX�&~�b� �L!��
E��	kO�mJ<���)��ŕ�9~2�OǱG���.����\VH�{	�[��]hd����1�Jh��
i�&z�
�2yf2N�k6N>t,v0X�����f����#�~���a�K3Q��J̠T�vwb�P�;�0ٌ�.��'9g�1�F[qXm�p#sT�fcBzt���4
���T>C� �,?��g�|3�(�Z����n�|0��(�Xt��y!�#�B�w�t"(��Aל]�/�X�)���{?�W�Ɨ
=өP��NO�B���B��Ә�֑��t�-l,�SV$y�BXg�?2�ׅ�����;�#C����w�ϋ� ��2�h�f!6秸��Q�~��]��v�p*��2��64^,�Z�y�'�"_��7���h��!'q��=��(�{��A>`d䊅�T>_��=��wQ>wo���>a�]�*Z��-,�W�ތ���g����O=~�B��pDh���� 8�2:܏����
vw���h�Ã��ǻ��o"\i@:q�|�lT �9�SrK��;��O@�N�OG��j$�&�'J��ɠ�Z��,�:���t���.��S���u���kn�����T��(�8w���)v���V�ׅ�i�\5E����߈����8����l@�GtZ��&J���G�K�~�+?C<��0j�C� �)#D�e�M�$+X�j�A@���R;W��L`�"<\��Ԩ��\=X�O�Y��'���꭫��Vik0�����H|��wŹ�+(�*tD��B��ymk'~��ߊw�cx�8��P��C7x8�X��z����{�cxY{�ފ潫x&����ڈ��~��v�8�S3���'�O����x؋��L���ݡ|\��
�IW35&b��b|����g>�p�}h9���k�A� 4�,�a7N>w<~����/~$~������h�\���7�ŕ7�F���)��(�)-2C�e�{?+�0��~^Z�::"�I^��nz"�8q�B<��S��| ���6��O}8>����}�^��;�K��p��C����:s:�I���0�Vct���T�h��9��GW���������S��ӏ���+[]�^��@xO��L�A�� �&~�b�K��x����tE�ߏ����y�Fߝ��n�S�V<�Du'�
\gN��{�<��Q�;���t�ų�OTK��$4�������(,GE�J��:�pv������N����Qr䰛����(����O�xXy���CK���2M�v6J9�P#2�0��
g���S0�Բ,��yR ��x>~d	Ņ��9�wʃ����`|��q$��Y�0n�q��3�;�/0�s��8�'8��\�y�a��-�Kf{�h�1��IiU�9Je(����ěψs�W.B*<"_�x ��'�j& ȡU�f1�+��/����߿�kW�:(����?&���)ǋ�v�����������
š�n}�B���K�� �����;p��r-�//4�x-(�z=�VVr���rjL�C�\y��ۤm5V���//G�,WoBie���#_BK�����Q��@ޘZ��9�N�Q�CDN�&�PFu��u��p��I���r����WC[��q���vA����㕯��FΧ��cy},��a+��������+����U;�5�����g�ر:>�;3l��1�������Xmę�J<|�x�T|�}�܉Z��(��U�7��`�X�\C���Y��'V�Q.K1��ʍ�q��nL/�������3O�1���_�m�n.�]���o��݃��9+��瓤���s	�>���8~j>nݻ�ߎ��ӌ������.�1��ZAH^:��y����g��3g�ŕ�_�b��;�l��Ȃ���ƙ����=��矉���� 
�'�ŉS�'N�{�9���آ_?��'�/���'�{"ί.ǉ��X]]�+W��7��mH��[��A��V2(�
�ZvsZ�Õ�� �[
y�����%A��my�G��|��'��N��(���3�a@����x�]�g>��x��>��'�3�P|����}����$?�.�Ӕ�l��]��O??������[q�N��c&f� i��3����Hq|a6?6��a\�y;n�ً�k[:{q�ڊ��v��%?Bo��?�=z6�kpC�0��&|x ����T>S��؅rح�Q�u��N�,�[�7S(�������Z?Zp�s>sŜO~@2��e�r^I�'@^E�����g>��.T �1���*yRŔB�x�Ʋ#���s� �L�e�&~&�ڣ�G�!��k=�BLe��m�8�}��J	"�����z��Yf^�~���ש�Q!��������-c͑��8�G����La��_>��K���[��E4N��(q��>�>�N�na
�<�ʯ~�7v��.ߍ]��W���Z���X��Q�W��ǿ��G�>�D� Ԭ��|�m�� �nz;S��p
��!�|g?�(���%&+e<�SQ�YB��Ō�(,��i4u/���X�:_���L����z.�Ҥ<l�@X#��V�@�iDl�����8�̃7�i�
�E*�bw8���i;�B�Z��}5�s���.2M����--����}{{'���+��v��R�8F�����2��$��D� S�^����G�Y�c(��}�R<���X'7�׀��KM�B�A��~:��{��?�1�����ZG�b��x&�o#`v��8��P�y�X�=�H{N�7�Bm��b|�����S��d&c�2�c��������?�z�l�cb��J��3��y<zf.���Z����0*�^%�AxŤq>���s�̉x��i�'cf~6������t���6�"����u��=����ql�B��x��\��3�ѧ�g�K���z|�=��M=˔+�
�I��_��|�K�@!8�VC1��@�*������.�^�
�e)�ht&=��@;��У�S�<?|1VPjeh��������c�ⓟ~w�����t2>ra)�sn9>pv)�f1������̅S�عS���S���H���Z7�}mo�;�%_�����A/�ڈSs�8N����x��n\_?�N�O����ƣ�W�ژ�6m;�T<��E��X���6h'n\oFw[�z2f�'buEo�Xp�%?���Ժ��3���ΑU1t��×�� ��0Xv�9�V�c���N��`(9��*���BN"W�,����"�i��������,#o�</
~/�b����%�ye�
�,BA�@�YXLj�Y�;A؋b��7���$�e\AK��]#E��q�P�P:q^O&��Lj����QBZ/i}F�- ��	��/)�6�g��c�Uo�0�g��?�a#�2����|-�͂}@���SxB&���>Ru�J7���qB�Fݕ+Ϝ��gO/�)�k�`d�h�K�+�u���D��	��q��>��e	��-�B�K颹������q�{��i�Fi.-v5��q %�)"M|�Ѽ�P@�:�G{d��;;TW��WW�m�sQ3�!h�1`����C.��(!�������^����x����i�%L��"����������7�Z|���9P�WNz1qH�0�T��.°l�ßw%R|6U�Z�0�4�a��_��ƣ'V��'�������斗b��G�`Qؿ��n�*�8���S'���]�?v>�Q���|�����F��5�q�ӊ���`:�(���!��G������wy#FN�c�|�#�������O4>��'�6W�+3/�9��,Ξ=����]z8�y�$���M'��X��8�lT�����w�;Ͽ˳�q�Li���ƺr	qu2��13�"}t��R\:��q�l��'��g"��ԥX���m�L�ދ��9Ӌqy���OTs�-�-�Y��ҩ�xJ��Q%�W�t���|!�@!)�H#���Mm��\��=��d��f�r�8]�Ju�Қ�c��8�P>F_�]��e��9��� +S&�T!���j�2��
�v��;�ӟ��^�.��l%έ4≋K��3���{4�y�8}�tLV����n�m��f���v����դz.xA��!�\�F4�%n��w�p�g���S��OJ"�]z�6�h����Ӽ�r���7XN>"V��;d��`S�֛��3�:���ʦ
q�IA�am0�'ԡ̓dR	�9Q�˼\{F%������vi�����G�U�ҶK��K��PEa��h�^]!�ߩ��Rf�y� �Q�����H��G�l���#����2=�ui��L�gC?.dO̸�ő�p�^�̱m;K	-��n˵�_x�R<r~%�;�*�rz]/����m��
��r��H��ɡ�IW��.o,s�Ϭ�'Ú�>t/�v��am�|���C�Q��������
�>�/�}�.�^aa�禄P�8,�V��@8f/���B!%B���>b��=,4�X�ӱӫ�Ξ>�.�Kϧ}ؤ������v��MЕk7bmg3i�!�n�l�0�çO��~����O~8;ҡ��F?�&�5�h�۟t �}�g��s�*�{q��Vl���V�Y,��>v*�}K��2�	~��`������k[qks+_�ўE��Q>�zω���<�|�B�;{�F�o^�7��{A�c�.O���Fl`�:I���v�������x���s�v��?<?�ܩ�䇰��;��R\ <��?�%��p������g~�g�c��d���>�W�l*��ٹhbeߺ�o߸/��j|��W��7�FQ��x��e����Eڍ�����߄�~/�.�P�H
�>��bA eN���o7ۇ�{]o�,�hV�2�$z����l��l�J�r*,��{��
4���J
���EgW1Rm���`Yߌ�w�P�W���[����ɅG�T�Vqe{�I2�&܃����P�V$��9��G?yb&�s��ġ�GO���<u:>��������O<�>v)�|<��}0͸vg#n�ߎ�݈��Z��]a0Q��\�U`<΅p���#'�U�@!e����
A)r<�8�s���l6��(0��ҘGA0��n�)��#<@���;��Ү��
��s�Q���I��*��6b��Hq)���rm'ǑBL�	�a�F΋S�l���;t�Fg�2@��9�h;�6>�`-BqM�y��ǩ|�۞<�����#�E���QEU�_$��L��Aa�� �v~�iQN�#Qa|F�0�à�P��²��|qL#�,��x+�ӏ����慷P�
74��5}�Ue���-���&���A������iz�����݊�o! �]���{Q��r���+�f�<�V+�A{�A��G�@AP|N���̡b��)(
�p�0-{��M	�!7_t��U,͕�i�$V���SqEB鱷�ːX����*�6w��+Wފk�k��f���X��!R_k��ʤ�-:���Y��t-�Kk���h�5���n׫1��Ǩ6�Ym���x��J<|�x�;��ܹ���Jŉ�J���R�����ݵ��%��>g��ɳ+��C��ز�Al�ݏw�Fg�~\X��'�u*~��s��3X�(�����׾�����|-���QTws���⧁�ً������/!����%ɩ8G�T�G���񒇓�9�[�,/����(����Qq�8����x��+��7bcw'^��z����{�Є����݋�k�q{���Q?��es����������-��;���9�|�ˡ�{���� �`�4�H*Qc�Jc�홚r�*K"Ȗ]���*W�mUy,�V�3$� �AA�@h4:���ݜ�=9��u�림�]w������+�����/����n�?�	��٥M�c�A
Q<	��Av \�ԝ�ND҅>�P<p߳������§�Ê��[���B\R�P��see��|���_~�~߾���wT�]J� ��㵠��ߨ����İ�:�ޯ[��e��c��}(w��.%�oi��Ϝ.ۧ�̠]C�і-����){��cv�䒥�Ӷ�۷�-�����{��i��
��g�(PU�nA}5#S\K��w��W��,�S��yC}*4N��)��G� 3TB����&BW��[���u&J�ݑ�\`��yF?q9Ɖ�T.7�eYh��{�!�>��~Jr��2��V�n)�O�� j����WYF0�-4���p),N
�vꈎ˨G�qY@�N=P��axI@z��r�\K�����I� ce�w�A���:�ٛ�g���pzV��p��/�����p������t)5��5.Ӹ��b�����Z�o_ߴ�r�"G �̩�}��0�;�P�,�2	c0kucG����^�����H<�e�F�Yʕp�����hup��M;�����Ky˕�0�%�l�+���&��!b B�@��"�>z��H&Z�d�~�
��LQ�����yK�*YJ�%�i		Ŕԭ�5Z�A�Į�������6�ҬS��-"W@��memǾ������!�{j�"sE_�����S����C�t�|���$S�Y;�P����{6M{,3VD��:�X�J��V*x��K6�~�ik�C��5L%�mZbԄ1n��������i�X)�7�[��Qj������?~�z�w��Z�z���v����u[CH�B�X�6�ܞ]��q�L��ʆ-�]��_���c%;h�(�fVm}o��h+�#�`�3%���/�`��Xߵ�^�m;{��װ�u`�&X}:�íh�(����L֞>Y�S�yx�p!n۵�}��ط���}�i�߱*���3�vbq���![�\�?���d��� )c���i��v�C�L��!lC����RL5��F��)[�aw��vwl�4
���ʽ���޲?��7��w�c)�-�>�lcg�޾���g�AK(�+/	ʠ;7�6��o�=����]��Ú��"I��q�:��J�.Kٸ�<�g���ю�.E���);sf�N���Z�����.�c4�b��m��g�ZӶj��R��>t��hŔe
	+��$
�Q����c�+M�"�4D��#x���((rM�s����C��U:�[��,ˀ�����]��)��D�7��K��	��,� pV��g�����8�,��[;�>����h[i+*�E��ӗS�)Y,�'Q�L����Ix��Լ���Ż:��X�a�X�(&�� ��2�uw��(��y�Sbc��g}O���^/�#&�^�������E�!���������ػ�8�	�k����
P�1R/'n\O?�4��H�;��p�~�?���ذ�3�'�K��������Ρ�zN�EF�V�jq���G�Z�6I;mZ��mh�����.�MSRe�T-�v���mw�m�.[1�D��%+-]D��I�߅)����Y5�Kp�L���E>��[;8	�^G����E
��.i5�׀��mm#�Ƨh�;�Rh��&��c	6p-ʥ3�ֱ.��M����mW����۹S�v��i;��#��#�'��o�_���f�0ҹ�E�S6;1S��}�eh���=EZO��l)fS������<�H�^f����r$HZ$W�.V���-�L�Ɲ���S��M��I��A�n����x��h�ౠ��&�ۂ�E���vk$n��������,�;L���z�{=k�-S\���/�O�䧬�V��+k�W�����_|¾��O����-���0�+��԰)<E� Xh����}���|�kݿ�P��Ə����aE�yP��b��}b�~�����~�Ef�����v��]{��{v��={�`��Z&�}�{�KO���:V���֍;֨�mvv����T*�4ȊQ���E9�
h�(Qx�K(�,�Rd�欅��j4�hkۻ������OY�4k�_�,��v�q3����k�>kΝ�Z�m�?�k�贕��!f��lɎ�6M�X���]��N�o��ljrD�)�>����>���s����/<fϟ�vfX�j+�ʎ����ڭ�޹L ��;[;��o�cVVm{�i�|w�6ޫ %�(L(D'�v�`ۉ��5�:����]�fZ��D����l���M����un��Y�pSsq�>3k�c3����t8%���u+FxN�'����)4ﴬ���+ϲ�\�d�����'Q���"����M_Q�!g��	2I�g�cDPL�HV�1��t:Cx_P�|�R��C�z�<y��g�Π`i��w� �,���λ��Tg�2����0ʁ0�Kx�֘�'\��q!L]�G�C�@�%$����q�b�JO��_�>VOS2��$�c�<G�Q�=B��V�Ƣ���5�����z3&x >�W�����������߭��K6�����/>u�N�D���X q������� ��9��ٱzmךXQ�쌕 j���F@^�����pQ:�ƥE�}�j�4H�V��4�۬���Qw?�Y�����|��	$�R`�`�����W,�x
����Q���-G�,���Fpʩ�4���Q�h�jVot�����kjf0* P��.[��j�����ʞ6����6� M�	�S�Y�'����R�ŋ���c�ԩ�.�f�f}sSzǴ����(����2D����]{��-�v3Y���gl�`�n-ߴ���j�o�a�Ú���&��:Lqc��Pi X���{�&l���ᚲ[��v��M۬��ZIX�!������N����Z��k���Kv�����4u]փ�؉c�fH�l�Y!��B6k�B�����]ۺux�E�Y�һ��U��͠�W��?�?��o����w�����Û֩��l�*ߴ��v�������>���Mڙv���+h�@�iLc9c����Ww�@����GYדq����U�:��=�ᑭ`�ܺ|���>�����.Ĩ�"o߳�~�#�J��_�c��>���޵�~p�~��n+��v����p?��j|y�>��m��vm�Y�����"ۇ6�O}o�4��[�d���'��S/<k3�6]��\n:���Ղ�l��HiE���d����]G���kM�mba�(���)i�N>mu�j�ЖFڔ���%��([��Ēo@WM��f�j��C-2��c�e��5�I�L-�+�/����}L�]z� .`�7�b�GYXB>���T��Š�*{݃���3_��~䣬\�p��,h�7���\z�oKA#�8�;]JC�4+F������y>�mu���Y��٢���A����'u����?~WH]�yp�����Q�4[��`���xy��㉃��>�OJ�� �q��L[-�M�2%�	�ew��}R ��,R��QL�ſx�L�߾�i�[��"ӥ��������Adqh�y�xZ8�[��uUq�Q��=��}��',U\��h�|�)PL]��Q�2��#�)�Ta����m�h��0U$�!髆����! �	L�g*��?�UD���D]ia�R�-?l��B0OKȋd�i�<.�H�I[L��}�b�*{�zdJ��sb�3�j�j�ݪ�\�m?|����[�2uJ���A�w&@�ڀ�k2E�Z���%�7-�i�Ř}��S��3g���%����"�y
�]�uΊ��j�i�� @�ȳ�����m��ܷ����4��ӏ���ϟA+���ƺe��z��~�k҃=m��CK^GN*/|Q��,��Ҕ6궿v߆�H�RQA�C|�3i������a�0����1�]:�E�$-5��i'i�����]ĺ��e"$Vװ��8�"dFç�:�[a�E*�#{�����-�w���ݼ��7� )�Ї��P�F%�i��A��ՎEV����t�2��@�2X�����*"2)JzNI�	�fLI��Z�Ǐ��0���>>4� W�)�1��i[�c0���y���5u���s�iƭQ����~�f7�V�ڇ��|}�YgF��i�X�#GHWA�4,/u���P���|�.<v��``p�����X�C�PU]i�F�m����뗯�,��F�6��h�!��.&Pr\ P�Ӗ9��5� j��]`�I�j]?K9�Æ`����!8N9�����\��Pf�YAVV�`/�Vyy��w 8z�� +�6�i�k��]H?�q�_��'��q��T"
���^�?x\)� �O팧v^Q�����7O#�<$|�,Nb*�JO�3h�/��s� �l9] "HC]`�p�2(M}�1\��W?H}�D��%L��å�`�ӫ���p&�(O��O��Y��=]��\���R	����()���%��UoO}$�!��)>����m�>W�[�.�4��Si���O�KO��20`YS�G�X�v��j�H��h���\��rT� z�`�Z�E��tw76-9��4n-�L�����}� ,!��MŖƢj���
7�~ja�מl)�XTbr��+��H��.��L���O\ ]���|��V����w�W������<�ZSoTm�����ӷ?�?����jw�aī��4�SGShZ���TE�@���C�i�lKV[v�d�ʥ;w�V��T�0���������%��l� �ew��>X���U���=v��������3	+��lzv�����}w�ٹy������4��f\���b0=U�|��*�ei�P��Q[<��i-<��=8���3��l��Y�@;x;J�jUHX�;�=�a(-HL��W����VU�P �>xGA����% D�"�v�:��m���N�Ѵ| g3I/X��I�y�1+�:G%��<MYzT���"�	����,I�o��D�j΄�D��| �Zֿ.�'���l֠���`�=�j��Т8�0.G�) 0�}��g�N<G��X'�
FR��pe��^��D(���Q���P`��|��\"i����\��� 9V��?6o'f��cɩ���D/jY|T.�E��n����C�������{|>�>nh� �4ޙ�X��B��b�7���1��;
��c���+kX>U�R�3��%`w������h.|�V�<����L�~��{��xS��p�R#I�zRt0�Ƙ���G��2jc��h��F�|�Zh���!LX K�+{��1�t�t�1qj���P��g����]��Q3�TF?j��ZG�޼f�o"���=M���i�&u���o�P�[�Ky� �P|/��OePq=wGO��<����['JCI�_������Z�R}tI�)�p���)��t���(	9��Gz9�D">��R�J�X��u~����>ژrt��Č=n�J٤#�o��f&��4�H�S#�/B��`q� "�J��+��� ��>�(��5lc힇��r$��s	���>��!D�|֔V�,r�K�R�����M.��:B�>��g����.�/�
�� �e��o�� ?Y9�=Am�cM@\֏�'Mv/���j׮^���t�v:S�;k���o��i/�VΒg&��E��Gh�݃:̶��'� �[��s���əiK�aP4�w���lyy�v67��b�;�����s��=����؃�}��ڲ"b��+�<GvX������V�����ʙ�=o3�SB��Zu}hV��8�ig ґv��_��0���#��I�W�̩�n���k��s������	��!�C��?Vm���+��u��vk�v��U�Ώ��j���I;=�h;��z�FZ��ɭ�cm�=��4"�5n&��ل���?�h_��S���>m�?s�Ν=m]�j�ns�tJ$Kz(*I��`��3:A�G����ұ��b4
1���)nM�좾o�ۨQǞַ)��^
�q���"�Gǧ,��^�M�Uc,
����{)p�;�90�`R�b��'܇S0W���\�.��-�$ ,.�%Sb���M\uv��`��ݹmW?|׮^�j޸k�ܺg+���!�TCd��9{��R	eG�p���تA��p0�*`B�Ne-5U����d u���<���ܫ�Op{��l�.�,Kg����'���_�Z�0�M��ܢ��1[ثSÙ��u6����b��w,��L§��z�"�JKm��\z�cx�3������BLX�����x�v��Ɗ�r'Pړ���+��e�m��[�|Һ����h�X|� ���xڡ�!/�B�%��W}�a��{s���*��NV�`���t�A=��ʃ<]�\Tm=��h{5��*�����䟒����A�),��o"|0����a�3t챴����,"�p��D�N�p�H5�0s�Ҡ^*!H0�[�v��,����i�]����Ҏ��!|?��	�iVRN�T2L��p���w{�0JG�A�#��7�M��.1#�*-��T���l���� x��C@wf����@ig�^\Z�T&oW>��Ο<f��9a/�I{
������w^'�� d��w���8@j>k�Ј:�0�梶0���8�Ս�XWw���}��ە+���ͻv��}{�+����ٵn����`��l�a�YK���%��
�ϑkAZ�/�Ѣ]�:��a��)C��p�m1��e��ff�,_��:Fǖ��H2mC�r�"��FoG`�U���+֢�)��,�]9�����
���w�ls���}�q�}����~h������'۹r���V���-<��YL�b���L;1�{4�0N�k`3��G��rjgTHK���Ĺ��rq��85kS0��³��>���$�O�Ɓ��-����f=|�\�A�%A����� ��u%ڥ}m}ÚX�bV���)���X� +f����5#a.�Bt t�V<SQу��8�*�23/G�$�G���*=��'Ogl���>mr����|�V��6m}}�sǮ]~�n^y�6�߰��-[on�[ǚoa�Bm�N�(A!�����"Ac�(X]����3*( �)%�S,w�O:jJ�mS��#�em�c�^V��	'�#�H0<Uo�9�%���.�ˏ�r�$�Mx�O�~T�G�f�I�E��sc��ko�p�u,�����.z��� ��:��Z����t� �@�Kœ�w/B����τp�;p�P��?8n�(�,�pMg$]�(�����8e��z���,�\��z��Ke��*��\�V�9�0:���*�_x���l�¥:K��&��묿1��_��[%z�{$A�
;����&��+8�#�������§q���7�����|�=~r��<6wr���VX6���Вh~�T�N}ͦ�-#0�֬#Ժ42�u�(tC��"o�I#h͂�����n-��"?5^آ[u�7��W��ߑD��qC�%��F���vK�B�&���)I��+�'�?���$��i_7���<�����y�Ο>nO\8c�<q�t�����}�O�ICIE_"���J	����i���y��E�ʨ3�d|d'��'b76v0�pw��߿l���ݾ��s��ulS�E޼g;X:��-;h�2�G�J���;uҦf`�,��s�����:���g�9u�D2-���F��Jc-5���(	w7��a�$ȗ"(�a����aD�6W�ٳg(C����*[^F��y��/߳�wn���C�nذ[�f�g�����h�iK',&x�H������˒3��d݅p�g,%qG��=~b�^E8�*r�ʈ��n�67��XFBLV�f8����'���.�1���?�%��z����#��k~���\t�k�v�[+I�9��	״�R��Kд��ST�!?l�u�c�P:~A�����ս{���/*ō�x�/�,�@��s9�����Ҕ:-�����oc��l���k�z�!�<ڷĠi�Ɯ���D��~}	�p�eaڇ-������t4Gk@��|Uhk&F�uŒ1_�+ᓛ��f5�z�e\�~f�-�`Oٓ%��H���R�4f�QW�T��ƌu	�ѡ.1}�s{��5�M^����O��V7o�}%c���f�y�F�Z�CX�#	����R��o`�r�2Q8�/1���Ixr�ْ��������n��S�R��3�O�Z/��<�%K �b����!��^J���T��>�G�zSV^z2U�B�=O���//�?�v���
���һ���uʵ�Xх'�����
�	ȃ�I��~����!��������੄��1��d*�ܿ���il�'���P$����"@C��Qw����5Ȯ����V�2�����\F 	!t��
(! KEw]*��êr��U�|a���n� �Fh�}k���4h
Q���4֦�Zٮ5B���%K@}���R�9��6��x�~�Ӱ�;mK'��87m]궷_��C�J��/ |m�/�n�H$�N>u�Da��Vd�s��!���{��1��_���w��W���W���/��sO����K�+��%���E��h������IW���
!4aC��^Z�$���hYC�?OI+�#Y�S�C�ڈU��em踂�t�:��իU{��M�}j�f���N�$PR��t�M�P�Iwm:5��B�f�c6��������r��m��>�4Zi?�Hi�퀫xBƜ�E`X n:	W�E�WrC �8���z�a�v����I���)�,���?�8o"ڱs��{��:ޭ�]x(�|��vOB��b�2mx��.�Dϓ`��W�~wx���2��'Mu=��Jn��n��}���? N�h��m�d���JM��xq�����|R���
	�7t���N�X�I����[@8�R����0����O��2�<P�1Gg����.&��A)�	��k�Cp��T���[�v�\X�5�H�SJ�ĝ4�.c��l���]"���}�^~?D�*���嫶<Z�]<c��3)]@�����~����R!�cH�_��~a����s�9	őO��d���{�q�>9ub)k��l4��枲Nᄵ��-�p��=M EB�#�g��"���SZ�C����5!ُ�q��W��P|�s���	�� �`Z�������=O^�p*��RT_d������X�A�s{�¢}�x�.��u����v��ܛ�#�!ڱf��+��nP��g��i�h���!L�Ym���u8�: ��1�D}�>��%;.0��0�#��(=4NW@Vu�i�Pݕ��#�� �(O�rn>�܂#=�Ir��Խ;��똚7�޵+k6;7k'ϟ�\)gG��ݚ-�n�;�}=4�h��Y°5�U�F$�D�g{���q��Ȧ��v���=��Y{���Kf`�][�+��O^�.��Қ���c���o�o�vApkƠ�Z'�.�M�dm_3�*%*!&�i�c5-��8B	�T�>y��&0�KKf���&�D}Q��w`���%+��L�2H�z�s��pk�SgO�+�=m�K��<�G��q:� cԘ���kZ����ރ#;ܤ=3f�Xa��4y嗥�I�[�Aʡ��TM����n��t��ϕ��E,�2����Xmw����ֶMcm���e��q<�;.�T�G�F�.��L^|6��k�0$�ǧ�_;`Ϝ<n���������s�g����g�-s��U#�֯��k�l�EN=m��O�����
СE�#;����g>a_���|�.}�Y+]��م��j=8��bu}��hL#����/=�dN�!Dt�-
	
@F�}f2��\�$�I4�1E�AI�`��Z���p�kz{���,�U95>��̴Y(zeA��j���z�B�4�e�IK`)��5�nA���u[���ָ妰���֜N�����7�������|U�����}�I������IIϔ�Ćy�?�>����E��L�9=�� �[�W�!-1#'O|>*A��'!�� ^~Rv�Ђ���ז=>�[8$�M�"��P.ת����J{��믺����zMyW����|Ŀ&�>J���m�/i�G|Wu��^����HahmNс�
�yQf�{T�Cb�8vn2��s9������k;����k�V�W���vn>e/������%%� b2"�dvʻ��[��c��OM�c�vz���<�h����b���6��塱��iS�җ�)�IkM�Q�Xm^[���5)�#�~w1� @�n�����k��Jx	1d��u���.u��]� ��&��%��j���oI���mX�[�1��-;�����&ae�"?��a����݊��!�ɶz�Q��z���O/M�����gW�߶Ã�E�]8}��g��v�Ʋݻ�N]4�Y}U88����<�'�@<�Y�Q��v��*���@��3*$���G��nQ���/������v*�є�h��^���#���G֪�d���%{��6lʪG����G���ebiK���X�ُ��;���F&�w�1�G�rON�ݧ�b,��'�W��qPC/�tf�l��G)�r&
g��[�vg�GMKE%����B�REx��BNx!$ ��X�C���e��-�:mO���}����_����^x�>��3v��9�*t�GX�<g��U��_����/�M��Ͻj_���W^���۹�3v�؂��u���~�>��W�+�����)��M�K8:,#�M�؆��pO�u<o��8�;dX�e�&�&eJЎǸ4�'� �:J�9[���T���OY��m/�_�&(:yT��
9�h̏3��t��[��f����3���nM��>��٩�`�����Y
�4@�i\yD�8.7��Vߜ��D=�uˏ�n��_D���Uu͋�k뢮��re�'���w�r��%��n]���d�n{g�c��������&���Up��&��x�������4T|��WD�+�;�Y��O*�So�#�##�U��?|!~�@��B�?N�JSah�3��W��O�"��d� �m�g������KR.|$|�$ �@81[Vֹ����7����mV:�?���Nإ����\�.���QdB�7�������)� C�o7�`�*
#L$���2]k��Zu-�D��QH����b)D��lg{�>��C��[�sǶ6׭���n9h*�	���C����㠾���I��ql/�����^5�N3�8��::Y��J��Q��$ԃ�2�u�q5nRG�=�4�+j~�h�r�ˤ~~m)�wP�7�䏩�r\B��ڨ�$�Ԥ�$h�=��w�.:By�Y��A�{��;���������{�]��_�+��Z}��
X�Z,�����);ur	a3�@l��s�v��q�k�{���X5�NL�g�aP
�s��εI��(}��[�A�i�:��@`�];A��S�߮Q掝����y[X�������X<Z\�KE(��|��6l���x�oG�!3cq4t�v���9�.7!9 W�"��� +A���.�(�-��e��/�vݤ�;���������a6ius{��dq��E�fG��0��X��f��$)�wa���Ś��N���?�	{����"�����,�۝�ekA�O�;g_�韰_��'�KO,ڋg��'�.ڗ?q�^|�S�[����N-.�g_|Ξ8q��3I;^��±y�\Y�_ko��%B��kX@(8�Χ/N٥�S�����ɐ���E��ɏ
��qM����kޚ�F:cG}q�	fA2�v9��M�
w�������h�����$tH�~\�'>]p����ڂe�aV��=�lh�i�x�0��|�c$JE%��p����7y��>�'Ί��":Tbr(�T�8m/�"0z���.�7��|��oZr�����w�䜛(ܸ$��r�A��W�
�����4�&̪��J �F�R<)#��:�̃ T�P�")�����$!G���P� `���N���K_T\�����6�>���]i��c} _h*'	����y����O��w�p���l"|rލn)e��4�9��O�X�'�
�/���*�P� �	A5�3,��R�h4sV��ZB��zFцŴ}K�n�f�"=�-ʑ�p��� ����,o޾k�^�i���uwݮ_������.aJ5�VG��B\��	�g	)1Q}��|�U��7��(�N�`��AT_��P�trEۜk���T�T*��/��:/���ku�V�mZ��oʢ5�ȁ���BāЦ�>~�AX��c���J6���AA(��[�b	+�������/��=�����cO؅���s/~µjKҐ�S��#���j!efg�2Ȱ���v!��\�ն}����>�e+0Y�C0Bi��N�o����ÖP�Q	��-+���j�}F�q&�� Nd"%���X|:|0�a!Խ�v�k�pK�.�B�CKã�60��j6�ցĚ��#uU{�@�^ޞ�()���!�G�%�0^����EX�A�	Pu�����j#���6�}ю���q
2v���.�:���v (�К�/P�|*��8-;>����30�0P7�������+v��VȒ/��W�A��Ze�=T��O�چG���9�n=h�^�L>N{�R((��R�Dn�Hp��]�T�����=y�N�ql!���`%?�P�iIp7��7m� Ҳ�>B��nH��VY~�;�y��.ćĄul���tJ��]A<M���{	�GÐ2U�"_�+X!��u������D��"A$0�4	Bx�o�A C�C�/tlx��Ʉ����qB7�W����K�^N��L ���\R�a��x�e!1ʢ:u��^EڪLk'���@�v�8j�-�c}�n�E��ň���M�:�9��gܻ�x��RVp8������*��G!twH��!?-2�tkQ��0l�/Rd�Fb*�>�@uuV� #Ҙ����RQ��� �ɇ�s�Mc0Z'"-�_D-$ӗ�3hH�gN��0��ӫY���Lf���4}�' Q��4�4L��+�m
Ax陳v����ݸy�vv|�Rk$�']n�� ~���B���Ǩ���L�5�M)��,͵C������ۏ�}a+�$|�q��@�`��qM�>j؍���i��~��G6l`} ���L�ȭ�G�Cօ�� �Mj�y!kI�Im*չ-3%���:{��i��g_�s�κ5&�X9��69�~��I;yb��X}�V�+��?Yo��g�%4QN|[��]�խ�B���]Y~bHj��CC�9#�ԅ���̯��8Txi*�LX��F`�I�E���R j��L;������a��\��-���V��+�64pH�� ��U7Gcn0!>�#<U[5`T��m�=K�gN�]`�m��Ҁ�,bV�'�V���69�k|GG,������=Y_�g}꒟��s�k;�SEk7Z���}PF�����=�<#"����g^�O���A��=�v�C�l��`�=�O�Axi_6�X ��b0��=�ߴC�	g�#�Kx8�GȚv�h�蔆���h2H6m��ehWJ�PO.a�pd�I`��0�0�]�����L��ʄ��|��]�V����0(�����������)?�+�[�
��yw�0�@������3	���@~��B^uk��<:.�}����E݉'kK�	���U����,�m9Xb��O^>Q@wUH�@7�Nʕ-��*׸|�����x���6������6��X�p���M�4���z��<��
��������nx�a��E����i���PG:��靆���Ly�.�p�� ϰb�ذ���i+%h+(�x0 ���UlX۳��!B��9���	)�r��	Ͻ��5:�3IY���X�愭u1b �[$���N*�6Ǆ�AF�/ Pr�ӣ�$#�q���45u�B8�(�hHG;8�i���j�8���w7����7��wmcu�bXK��\�R��p�����>�\8	� r�X6k��< F ��@�!0*�V.Da(5;8\��с5��\�Ay�~t��Mӂ��f*iϕg�թX�O��h����t�i!�5�:�@Mg�o���sa.�����e�k˧�J�YIH{�1�R
�Ȫ�:�|�00��&UȒ�$�`eH�Vק6�J��tb�uK�*;�#�����y�	%�	|VY�!���i���%�>�>\����ّ����I�5����i��LK���8	u��n��-�%܁
N�Fk҂����4m�r`�;����o�;߾�h�.�_�{�?���˦E��_GL|�R�Ne�.\8gg�|���-������o�ٟ���W���@/��V`Ph��<��~=b��U�;��B`�/��R��T},���Ă%<e	�"�,��v�e���ڴ'�2�� �N]�}�?M)��1�.�w���E�;�� 4��&�M	Ͳ`��J����{}S��]Ci{{+���\!�4V�N܇X���K��U_�I�^����]��>,E�<��J�oP�y��	�#?1\(�����0q
,�I���s��9��a�f��D[��	p>�@B�Ki������V$��5��|U��]N����?��q=����.�	���/����`1��<���0�W�ه+���G�%�+�%Wu!�YG>V0�0���Z��D�����74�j ~���������V�\�DU ��H�QE�pKa��Y�#bl����qI�QSKs�b�{�bW�Bd�-�K������޾e	��v}C
��$� s�]�����)� P�#��	R�Q�b��71���0'�rɮh��UQYP}4�}����=���oٿ��v{u�r�/�ĊDSm��tE�,ʊu�r��C���Xan�DOk5�:�?jZ��n��5�ܫZm��´��ܓ����pڲ�i�o�����ح[��0��n��5QG �:VN�(w������i�6H�vw�|��k�J���L3Xhb.�R\�R���X��QR�� !���Gڸ@����{>���T��U��c��
����U�ߣx���mq� @�uJ_]��s�}̈a��S�A]��60|�h������ڃ.��A�8x ��9^�[B�x߿kF���)ߴ��&�\	0�X<����k�?�l��\���u����A���u���w����V�ݵ��C���f?X�k��������ط��V�Y�A�j�Rұ�{i[y��]{��H��w%����Ѓy�n ��n޳w6W}�K�D��nXKeAK9���-��v��|����,��R�ͣ겤M�"s8;Vy���.�vr����/�c�ͭo̵z��z��GB�a�;Ο��in|�g��qZ�:mR>����o���.��Aa�0E��~Z<(G*�a�7z$�u O�y��+�<;���4��~^UQ�|5�\*Ou�H�a���"� xD���4�
��GJ���^� xtWy���8פ�͇%�et�/�A�C���=�2斬�pB�s�����0������yrc�I�\��Ͼ���~���G��Y�'N���^<e��ZDH@+9E��d�,WБ�s����s��"��{6���ΞkJ.dp��w/��DTQ1�Z�4+@5�۬Z	��m�`�kX={����O=e��,UA�1
�M%��a�k�^a[���>3�|�D� ��P��쀤���Ob>ҚZ���Si�:q�~��U��{�{3b�٤���Z)1��m-}��Q�y`�����"���u���@Ϻh�Vm�in��{eЌʔi�D��n������k�[�ܲ��V���{v���C(ʂPU�
��N6��SW�@�W�#�$l:m��M)�PJ�q�n�;H��V�B�:]�e�T�5�
ƆmS0�iT�F�f;[�#b���<s�N..����*vH��� �����#%�V+k�{�݆֮@c�Oio`!ďaA��'�m5�Ij/URm�8��O�94ߥB�G`/��^��}-�=���]�!�ր�zԦ��B8-��v���Rf��Ѵ6q��k�����hb!9�=�!y�P��õU��ݱZ�e�_�����[��w�ok�޶�J�N�(�L)������|˾��Y��7�m��D�h��ƾ�o���=k#����-�?�f>�%K��s����5�n�W�n���<n'���Cp����0�vo�֧ve Q(닊u���ߴj7j��~K[=���
��E��6]�sY;B�Є��0aM�:@Rc?�aE+SD�kcQ<t,<eC���P"GX��Rʢ�i��n�c������Qw�/0WK;Y����=\���.��`�|"�4����nU�E!�|ޝ��g�;Q�`������)]��L�Eg�r\(�<o	���(�c��!�$[@g�a�"x���S��ixL� ��a���^R?�H�_U������n�o!�P%��/�D�I�
��7?��DF�&#��:|	��De��I�JLx�Rk�^���ٯ�� B���_��Vݞz*c_{�eyª ��Y.hX�G���������m��m�܁8+��%�_۶���PL�tPE��Sq�Qͤ�⸆���q2KB�to��F�;nO<��=��V�_��*._#A!!D:<�
tҖ��GoK� u	%}����6���\!+ALGi	���h|�H��k���.�,[:osh��-��M��. ���!χ;���\����9e���E4��&W�X
n�Ժ��mmq�`�6!�&�C������#;QJډ��;q���e�ɜ�<>g������p�6v��V�o5تI�lvv
"O����򄽙��p���@0SSC4Dv���� ���L6� t�������'jEIKuw�z���:y�^|��,����u��X����a��R�F���q۫���+W���	�`�h�6�BJ��~I��[@�*����B�hR	�������0���d�F�;�5�}�C ���[L�/�!�'�����)��~w8.��-0	'Y�ꖕ0�Alwn`�^�fo�������{����}{��߲�;w|sM�}�zyϮ=ز�����{v�O�Ԯ\�f߿\�7W���Ƒ]_Y�[+����;��^��[vg�e�]+�2.��E��B{�UP�W,�Zq.c_y��-�M����m�_u	�N�Ҭ�?dŪѵ�BZ��*��v`��Z+b�-�\�0�eVGۗ2�@y�!���Ìꮯ��:�Uq2Mx��Ll�[MhN�q����S�t6��I[>����>��a���)==�0~g��e�Nc��n|
̑�B���2 ܁G�r�/+DL�q���},�q�R(������w�Ox��G�䚔Aw���?���2P��������/�W�՟�tjʬ���������z����|�}��]��	�1��b��U�&�GA%;�,X�5;��Z��'=w��9���� � ��u���C�_�k���_����rѷ�Q��S��\*E����rG�=��M�,�/ZX�jս}�� Ѵ]���P���K��g.�� �,����)�K�+M��ܢ]x�1����p�8Z�ab�-���)�4�|2�vH��-��1#M�i%dSp�b"���	}��e5)�z��f�#;V�Z:�`�3�v5R�{S'�wwծ];��U���v��`6�$0�Zl��x�B=���@���"�#tFh�q��]��=���l���lq�d%�І��98���d�o[[�`��]�~�h�xRC����5�mHͽ�(�(泖�J'�f��sf�lSG9����:y,�RY���������|vf�Ν>eO]<m�]<cg4i`h�;�F���ɓ���OY	�g��3�mjᢥJ3��>n1�c��l�d�xѮ/����͈`оb}M. /R	pF�@��V�s���Ț���Y3t4]��Uv����a��~�i��ح��mV�l=�Mj�<�5M@IF�w-i�n7v���R�B��V[�?�Kᑵ�{���A�8�T�2��RSD�F#��!��Ȏ��dn_���uTꈂ7Tиvx�fw�?��?:���޷��Z��۲���\�"Tע_M��o�T!�#��R�³��73�Z�[<3���hř9+��AGK��q%2(XE�ދ�6Jh�:7���NǢ]�θ���)jo7�M��BQ�qG�D��,��.y	�
IN�N��u��!x{�5�O�g�	�N�,Z,X�����z�ͻ��r&��'��s���"��K��ϔK�
*�.���6�C`�j�x��>X�q�	�V�ΘqzW.r�yFQ��|�%#��B=�g�t���[���i(/Aٕx�7Ы�o��C޽�N!$���s'��2�io9}��
&r���5.����؅��.���{9U�.��h��O� ��@	� �ׇ�
ϝyv˧h����ڪ��޸�mۗ/��/��L2G�Е%ȪBˈ�f�TH}��3[,��e��mGh8��U?����X�8�(xK|<�;�#'t91~1�"���[B��B�עF�  �P X<JGH/SPu��#/����_M&%�
�%?�v��?����?����0�u��w�ܲ;���Y�h���hv�U�ܧ��7�f�+�m�ջ�����G1m�X>�Ě����(µ%a��Z�f��<T�gxΕJVFx�����捻��w�?�b�~�m{��ڇ�g;[0l����<j.	�'����4�lɋ��=@J��f8�wf_k��Z��1��uu�y�k��|�-���I����1�X�mU4���4�c�S?�E�[�'��ӟ�ǟ��=��s����_��_z�^}�Y{���3��ک���KϓvƾׄQ�nR*�y���j��������GЖ`ئ��^���74+l�m!ԩ �S�P�e�X�I`5�8���hs��8�L�Wk��� *�b��n]���ޙ�|s-8V*>��i�qQ8'���J+���e�F�	�@���q�"y�#�/i!"�P#~1c����%�Q��WfP>�*�=o_��v��y;�}��Wp/�3��>aO?�=���ؓ���g(W�j�Ly�ٜ6�v�Mݪ�����QK�㾱h���(#Muv�ӵhC*��{Аe���x9��h�i����H�QKꀺi�Rٚ��K�jv�pPz>�&0G>���\��Op�g�u?�N�|�M]1�qR%�������F���8��R	��E�������p�k�����R۫Ԣ6��!\�"X**��o���K	�<���]�ht{ϟ�(��X�����TQ�'���u �.�%$+��M�»�S�Q/�A#��GJV�F	?e�p��⚤볭R�.icQ,�J�~�{���v��g3���O[ZL]{��U뻘�G��sh�+hܷ���b��5m(�P;���M-��R�Z�"B΢-�%p43���@����l�4i��h
NcK�/�#E #S�?AP%��>�X`��J�����k��~b\=�!����OZ��5�X��[B5��j!a�߱��������?����C��s6=}��z��-;{�EGV��}�\�N@t+�X]Z�_�U�pC�+`�07�Y��A ���E�7}2�f��T��/O��sWGS_�+�߰{��mgg˺�
�Ye��ō�"���M�,MO#��VG�iO-�_	�$x]�GARZ��X��5(F�V��J�1�� F�/RXnCH]7��«X����a��3��~�K���ҩIh'��r��)1�hWu��gm�<�*���U[~�mmڛ0#�nmd6J#l��f���!\���ԅۡ�Ҽ�5�B1�ރ�Fp���~�~[#�6���t�!5�W!�H;ިݥ�$@(�OLњ��W�(�݅q_��0�'<��{���Iw�G���:����.̂����'�C��X�E���GV��)���Z���@�jC�Em���h�f.������}�g^��_x�掝Cp�QO,9 -HPo���% @忭Y,��c�,Y�"����KDlg�a��q���E>�RVgԍ'��E��~$�	+zL`�j�'�E� L[�����Yl�kIʚӉ�R�JYk��
�ͧL��"�o��������vkp	R�
�CD�zV{Ji�q�|@�������Oa�4x�r�j��Y6�q�JZ���� �{Z��3d��
�v�.�e� �.->I0hr�'��"zt?r��f��GX�*G�i�P~�G�w�RY\9��O��|�"�~^?yA��>~>M���1�e�^Ǖ/Yt���-������<DD����H>�6��
��%K$\�J7&L$��4�?��Kg쩧_�O�j3�0�!�íu�Cz ���=4g�I䓆�t�L	iHZ�'�L`�� �A?zV���+��S*!���8C��ڃ�ma�T���_�1A2��h�J)�~H�����=�d 4E�5�;�m��ew�=���mۺ�f�tJ�����m�o���x���36�/X!_��l��� :��"�����L��9�r��xj�l�d��V|�˾������z�K��~�>�S�`����~�o����/��}�_���?m�yG���H�<��u��#�tM�P�[�r����Z>���-h'���H�l	=�y��К���T��νU���.۟~�M���Ahl���>1�����vn�@�a��%E�>kR��V4&;�R"�t:��qƧ�<h�ο*���m���"ޭI�H�!ȳ��9B��0G���nۢ[X7;�>���F���R��N6	�{�}<�R$s���x��q&�]WJBT�&p�Y]��MC�"Km�4��Q����W=��|"��-�L���YG+H���*����>�[�;
	t�MF��A�]���g`�)�:zb�����g���cv��q�W��Zb�(���3�x	��Y�Xr�E=���M���:$�������&U7���4���ߣg�QYh�.���L�;!���ؕ�Cz|W�y&�?���I�����gR&9�zp���sG:n�������3D�.-��$�;�*ѳ�a�yVJB�<*�ޔ�89]�ua	.	�nmq	6���+ާ8��V4��%=?:�Q�c}���rpxZ��)���3���^>�6�P\)_�j�+�Z������T:��y.�?- �}]c>0����-�6�^���<��+�lr)sNl�ȒOdK#A���ݷAghI44��/$U T����w�� -%����\��ǻ��,��ᩨ��r$%@��{gs�n^�lw�^���-��jvP�2��%���tC��e�H�u>�_傁��E9Ŕ�r�C{�UX6��Ʒ߰��M{��v��;j�J3�7,e�'d(�6U*��� ��Vך�m�.�)�\��♑oM?���{�jiϭ�5}�{TH�"�͟/�3O��|�)�_��W���߰_��/������~Ѿ�ʋ��Ͼl/>��]<s�N_��t&�Q9�$u8�V;W��J�Z�,m]��/��1��4���e�l6|���^w��sD:'�	�8������v����nZk�g:Et�ӲJ�g�k�X0`+P�y{��',�([���Q꒐e��X#Mڵg��=��|�޽yϮ-���ֆ?��pL[wC݁0~Mpж�u������On�<��kXT���ܵ��:�m�ġ���si�#�Of��G��(�i
ځ�{f$f !��p;�Q.����Âg]�v����:^=� $�����2�A�:&A��ݫ`>��#�HɆ10�Y�O5Gy1q�>77K�W���-%-���Ϟ*س�,���:eT����s�@�&���k��5Q�궶d��^�+��l�f���5%��X'���b�*�hl,�C�u��P�@�)W�����.Z��nC��h���!(t2��6G�n�dM&���X���D��K��K_�H�����]�p~�+�K0�AtNl�>����#�q���J�g�|�T$/��*=��{x܉�U�=����*��ܢ��������/�;���O�����5�u���tk}
EP��ƫ�j�>�SX����*�`���
פ�*��Ce�*:���D['y�h��&>/B��!��Ҏ��x���zа?x�>���~�c��S����@פ��|�@���X��7s���9@%@G"��S�]��a(h�=$	�)��3�߫F��n�hlG`S|ewϮ_�j����Պe2i�__�$\�ʾ��"�Er���Tڮb���F��&�B�t�*��������� k�!�|Ʀg�V(�!�."|���?��-N%����v���s,��7֎,�3L ���A��l����ER�i� �O��дb�(�-]Rv�Ң}�O�/|�s��W>e'�!`N���n���B!c�r�Ӝ.�1ۯ����5p/�-��Z�Q�O�����vj�I�$si���v-$�vlj�Ο>eY���E75U�oug�h[m�$l/&|VՀ��:L�~`��=��Bߚ�m���$G�{�ln[��G7���}�G������9���cs�M�m�n� |�4�I�B�D�O<]�D!n	,�!��E`�3ڤ>(�˝x��X=��@���0]v���,�uHL]������DCa,Q���_�]i��]��	+�i6>.V�`�a5�膑"��F{��V��C�
�F�'��M�.a�g4q��}Ɗ_�i����姗��m ��t�%)���\(�|�>Z#�W���SY�+Ĭ�X����"Ex#�#�kԬڠW�Jm���������=,������:D��(�N?L�;Zr�&4�e�P��jsQQ$�j�[z*���Y[��6�b�U¬�T&f�RڏSn���4a���`;��K*���v�6c��;O����\�����zX���5���xJ7�#}����gND���`��D�⋦�=��Rj:�6�1��BM^���`��d���A{�~�{#!�x������/�r됲���@��*հu��ԛ.r#��I�,?Q�C()���<J�h���G><�rn�MhJ�M���{��������'�wT����_���XFf7B���2��
0�639�X���$��T�Zӫ��we�ڝ�#� P�uR(�>�x��ƅ�(�V�������l�d�Bk�a���+��7ߴ+�e���������}��U{��c����)+.̑� 3��$\ �SLH���L֌<�_k��5{�Go����+M��RɦI���sv驳��:g�����>yq�^|����ſ��Z�p���G��n��v��-%���Xf^(Z7[�]��:Ikf����qv(#L$���Ϝ�_��W�g�'lj�`
��T�*��u�n5�Ta"��.eKvX��7��=����{V}��Ν9n�N�D��h*��Zwg�.|&*�u�<D��[�_9lՁU߲���p�NݚV��rV>��c�	�m���!u�< ����Y��g/����A�����l���O|� ��M�l�5�g퉩��_��J?k���=8��3T�����F��v�S��O�����}�ڲu�=�����u��1�Pv��:~Ζ.��KSE+@}�Wly�.8ٷ�y�\6��E!Qw��`�'͍Kx)�S|Aj��0�@i��Ӷ�[�M���4�
�������=Ӗ�<�h;wV�S]�x)������%�s�F5�g�`�>m_|�	�����cǬ�U���w����?"<�6ܤ�4`Adb>�AP��b	+<���r�>y*k3�I>9��T֒Y����&2h���1�=�bmcߏ���{`";m(�����&w�X�Xy6ag�N[�Č�#����� �7�k6v���36{�`�s��`��[W�m���Ҕ�<��SE��<n;ڬV������]�/8�0i���Xp���͹��;�o�Y���3U�˙�����/"|�Åo�4��sw�>�B]�g!��CW��7N��ym����G�{/��	��MB��ؓ�:/�Y�(E.���� shh�7��"�&y�Zb�>�z�S���J�HH��K�W��F�198$]l���<��21X:R\Yզz��y�4k���������o�.�_�������W|�hB�2p�K5
���C�[�f�V@��P"A��1�Y�u3L�2<7��HK�t���(T��7Ih5�)�<Ha�-��P�%��%������]y�M���I;��3v{�bo|�{��i��_����!Z����~:�EWKD�ц#V��øq��n�������������l����>�d����O�O��^�0g/<q�2�����߷t锽w��EV�h�;�F-e���B*N�W,�A/bU�d����[
f��oH}���}��%��?�����~���(�g�F�v���*4<'�ݵ����}������|ߺ�{6�]���i�-��7��l0~>�X毄�#�M3�X��ZEZ���t�=u���;��ʁ`s6��������G�|���@����V>9��!É�	R�iH�8o/=��=q���l�1@�OYa�l�������h�xoا� �T��>i��s����'m�%�㍪][Y�ͻ7�޽;�-�߸���8}ɾ���������¹Ǭ>��7�i��������m;u򔕴� kGݰ�q�����"uW7�,�i�@�~o-pPk�������ŋv��'����R�bӿ��[��t���z��c������'mja���*�0h�s%��X�<� ���F��].~�Ƚ]��뤭_�kN��Xv-�ڋZ�씽�Ң�9Y���Zfжt�e�h�ʹЪڢ��;�umk��6�5C���Y���`�Ò���X.m噄�97c��3��o�`�>��V�b�H34V���H� ����~�c����e���tҦN"|N!|b�hk��J�?�\0�����������M���ߘY:����K\��Qm���%剿�?���M��L�hB�&V��$i��?����$(B�]���Q]��1�i�@��2�]�Ww9UM�ԥ�r]`Gc0���I<��Hy��"�Cx���N�8�%JO�J_!��_�
'�Bpi򇄏������ڭa�;7 C>1�S�"��	~.
�eq�b����������o܃�v�瞝�g��0�<B��R��$���nݱn�B�����t�VA�hi���0x����h(�y}�~���- �-
�� ���� Hirנ��ƶݹ}��h�3�%��v�����=��Μ�g_|�
3��2I��-Dh����SL+Z$���ޱ#,��|���翄P���]�ճb��pH����_��䯾c�)�d������6B��5ʤ�K�I
¢~}��:�nGSU[�����8@�JG�ZcV��W���?��c�[_�Bj��}`�Y|}��;�����[o}`�w�ۇ>�� #W��&ߏj-k4;VCk�G�l�������4k��ډ_��2V����ê���	Aci��fln&gq��0Sl�\�p`M<i�N����{�]:{�>�ɗ��/�l�?��=�8~g���´M�-2(٬�`э�:���$`���a���,������ϟ�g�F�:_N�'at?�����O[��!��g^�d�'?e_�«�s6��}�]�XߴLF�s�� ۀ���H��F ��Q��U(�Iʐ�(0��i!�ۭ���.���Y,�O�K�.�b�hǗ�����ʚ��y{�����|�>��Y{r�d�y{r�dO/��xA�#��i�]6j�F������u���C��G��c�C���+(#u�z�ְ=p`�s}�b�n<�w?�o+v��2��X"O���~���&�x��ʒq���MO�-U�[Zo��ã���]={�Z:n���|�aM���FY$oMQ�pe,t���i3^?t-��I�e�S3���|���ӿSޱ��RlŃ�è&���b����_x&-���Q�Wb�e��t��$�_�<')*=w�Ç8��F��,��r�#�Ş�]e��\J�%�n��a*���2�T<7֥��!)�+_�G蒓0�G�UHC`��>"���������r�.s�?�λ������Td�M,jUB+���� ��QPx�3	��T@ʮ��,���A
_�%���12�&���R�C#�ᓷ����(ǥ��XiZ�v1�L��:�U�rD��� �I��)}���֠�6�u�=���`R�.\�d>�5p�$��F4����4��>{Y�k���ߵ��kT���N���ɋOYF��l���T�͡mo�E҅�4��[E贩��6m��ۨ֘�H����0Lw�x�4����T|�O9�V���[���wߴ��a����v�ڇv��f�O��m���F}��-�G �؃{[�&�h��%,�i�gg����la񌥳��<�mѢ�Kf�>`����>A#l3`/�!P�����c��܉W|K%M�� x������4��2c�Y_۔8�Fsm�c�<�Z�P�3�N��F����'�mna��CK'�v��1�~,���͔
և�ʄQ���
S�/Ѝh��4�jާ���\c/]��_��{�쩳��M��Br�t�!.@�A�P��h�Y���	��Pq�x4�O��s&���r�Jm��5���<id}��Z���"�S}���0��j�6�ŧ�Z���X�A˲�D��.0w����9�Ŭ�F�z��]���K��v�<k�T���xΖ��Ғg�ۈ���V\\��b�r)���SR/���@�����Q�㎒L`SR&LU5�w�U7��*`-ت.R8U�#\J"���1#�K�{"��� �\�c�q��M�~����H_�sa�qE	�M����!����O_U&�O!�ό$Ϳ�(���wŅ�����C��C(8��r�p�~A�y�2%��"pM�Kw/w(��I���|?�`S�r��C��Mq�&�6�.��k������$��$]<�w��|C�����K����E�k� �,�I�q)}��Q�ڕ+68܂�j(�2�!$�G �$U���Ih��HPw�v��Ѡki2�I�m�ڞmnj�в-ߺm+�o�VK��AYUXcb�0�Ũ5�U�v�����w!��=mG��왝Z<g_����B?9����nI�0��%����S]M��[0��\��\�+Z���X!����ҩ�:�!g[U�v���������8�V��6X�)�䥓L+��i�#�h���'g��Ỵ؄�6�k�	޶vж+7��Wl���tb`�9�A��t������lO�mh��C/5�*�C~Y�\��~������쥟�y+<��.=m�O=cϽ����O~����~�~��~�?mKǴR�h�h|Ξ�z���ۿe����������e���|h���-XH���߳)�4mK'
��c����.����z�֏�vg�fG-�0�M���w���Qٵ��]��}D��W��H��2�fl���i�X�`EqaP�LB(��"��mWĪ��๺;� !�r�����eJ�t& ��D���5����>�=�̫p��4����x�w���*u_W����J�)��ce� �ju�[�ZLڵ��z���C:c��x�z�]���0�-��ᨌ�e L�4#m�%!��fm����Ry� �i;���p���V���EkĀk�l�����±���6��L$�>K}��O&�� � �����_ʨ1_�K]��T��@)���OzO_��7��-��TH��O]�T��N�}�6g��)�3%����hY]n:y�ȇ�4R�5Hd�`�;>�K�0��qOR�Tv��Sr.,�s��K�Dƚ`���{����,	�}T��]�*Ѐ�(m2X�*��yW:�U(�J+�D����
_�G>�f��I�gKʻ+F�$�Ӆj&�𮛠'���KW�w~*���Tn0L�r`y݅���w�����g��P���='��/����Օ �E���
��8p�G�U�RNqaBd֭y� ���b�+|�U�-i�9/D�w( BV���4/}���pl�Ə���������k<��w���?��ݿ}���#G>��:iZ���h�(�����O<��}���_}�>����~���W_���9���t�%5�7*�lQ��V����)4��g.X�4meꖝ�B�'�`g���ѴS���W�v��*U���4���,�f����&�-'dv
��[����[`�	�S�'�^��d�э,EZi��A록�*^�[��&¦�z8�N����ј�v�M��	k('�Vvzvo�n�:D�H[�<m�Ϟ��O=e��Y���VoŬޡ���+.������/ګ��W����_�����[���y�~�g�j�^�,V�y
>e�^̮�D��~���[���-bM=yrў�x�r���!��<8��V�v}�b�{U�?j`����}�|��k�����B����[�d;0E|br4{M*�w���}�=�6� �>@���"%�rĽ6��Z+ZC>�.�Ld���%M�m:�U���:*(Zb�
;�B��$m��%.צm�7mo�K�`��{;8<��;-{��{��=��w�4��?$�J���6X@X��W>(1d�Cπ��Xyc�'�R��B��N���Og��MZ"�P�{݄�oFl�n���)�t�x���v~!kgf��%[���-�d4������'t�RL'�"LN#�@�}��q��O�S{�E�p�ݫ��g���.9U]���'�.�@BC4���yE�a�R�b�W(�M8�����m�iGJ~���7j�`I��w�!�.��(���#���+lA(��>)@e�)��ԎQ�3ܗ����˄�r:<�M��\�U�K4���Y~���J��..��Sc�P"�8�ݪ�Am5{���1�CH_^���x�s�S
��wb+`�Ο�!�RwsOJ��ה�i�)r4�`� `�	'hšr��u�V�_�g��ё�ٜ�|�p"y��g�D�Y�]��@a��0����Z�Y�YB�n���0�b��ү>\�;XZ9�".ف���u6����t��g;{�=��3��KO�cO<f3��q��hpM��f���ʴ���l��ζݾ{�Z0��{�>����'_~�>MZ�{\0�{7o�L>�Z�	��C�"<3�r���-Z�M(��+t��#�iG����1?:��V��8���n�D?�8=������{G}ۭ�(��j�9�]�k�w���1�A`��	lv�Jюem�``˛5ۯ��FK��H֚����
[{om�n�am,���?��k��?�������?m_�܋6C����P�����E��!�"�J��SDg�>�H��9>7m�>w��M�����ڮ-k',�V[;��2B�T����ch�|�u֖����b,��a��A�F�M_Ӌi[1:9m��L�{v��-[��l��pF�/�Dؾ�	jy{h?2��*�N$�ԉBD����Ă.���B�I`��|l-�͂1����۳��kQ|mUԳ͵U�k
vu���m{�w�o���/�m��7����^_;��V!$���@#je��p�Z�t��9�o�0+#�	����9_��Ҥ��Q٪�G�!�
i{�ܒ=uf��J&�FhTlr�7��Lka0
K����ٲ�OM�\v��)�km�&Z��Mk�daBC���*ϾK��[�"F%�"�Ƴ�$�?���B�)���
	%��Fѝp���˩��0�C_A�ت�4�MɏbU�@1������n�M;' d4CqD;
��5�>I�(���H��3k��#���^"d|=zR��\*ay�;N~�G��%�q�	�Tes��k$B�n�p�O����m��K�Q������>.(��8!��5��"c��~|g�ߣz�$	���RY���YZD�C��P�D��Q]$���u�����x�����l�uK����^8��q�ʞ�vm}�ݰT�`I���B�ݧ�P�#�U���C����O�\J}Ȥ��s^mΔ�Ƶ+vX�Zq�0J۽�w}���,Zx�pTn�G;#$�� DU?���txYb�Z"���#�>Qi#�������h�k;v��{x��ڳB>k�\�`��O�@�e��ܴ�{�!ʒ3�4y$�t�jM����|��T��4�!7}��ݷ/��^�"S���ì�h��$��EO�Ɲ�lƛ����aĚm�	�\�ٔ�����\ؠ5����m�8�����Q�*X�&PR!��q�ټ�j�ĲV��cxh1���"DsҔa]����vhh�/�=n?��9�{��E��W_��N���\	��2���=��rb��aº�`4rO�-.(�yh͕���Yݷ�zĎ/�/>J�������0���a���V%��[i ��7,�Ā�k�'���|�'K� �Vlss��?�o\�a�{�B��[��b��rv����o׾���[}�b�\���>YBS���|�c�V"�#�y��J������u�,͠�R����Z+��ٝ���{o�mo|�C;X�qv���Skb�mmPf�������-{��* i�`<�k��~�����;+X�XI �F�L�y��5ٍg���<B��E���-S6[J[�%�zP}��N�|1=��GP�x�#��Nmd�fʪ��a	�f	E!G1D�N�����%&m�ߍGײ���X����ֈ[���,��-^�[
\�`�i�A�T�*y�q�H���?��ӻ��&��g�9���R���Ԅ'u_�0�%�1+%���1�zF Ҟb��#�o���Ǎ9f���B����G�t���s�~�^�q&IP�lu���C��O`Q�%���'_y��2I���)]ޝ/�gTf��'�!'�כ+����c�7���z�z�����σ�SN���*cL=Hܡ���)Ro�AĔY���磋g�s(�N��P���?���6폾����l���~��Y;}|! ��֨l"x������mb���T��u3A+��
�E�.7�/�e�����$kn3�ԭV����׬0=e��_r+ek}��)+�W(�<�yxq�pB�hb`��c� jH!�WT�$o-��>a�ֻm�F;�z��}��UK `곅���?�v�	����Α�?\�
Xa��V_�I:�[{����cA��Y����i���]��-�s��z�SZ��"�c��P-Po�=��ð)�nBi�:L,�w0����sV���F$k�Q�6x�Csj��t�FV���S�2�ό�`�b^C��mS0rA���}���A����]Z�b�Ђ#[sn�xI�(q��{��l��
�G,f��i�6�x�B.am`�J��cy�;@p����B�Dq�u��v,;���N�a3�Na�b:Z{��z�g�
ӪZki�SAtNbԶF�ao�w�������7~d���������oٽ�l���[XWW���������c���-[_���G˧4��'4q��w���'֔pYkit�أ ׶�6Ee�ހL:�b!x��+��+7w��x��웯�w>?�k���I�G����fwQ|>��m7�sۮ�|`oPN�B�����v��m���>���#��5���VD���5��(mM�3u�F�g$HSvD;];��N4g�l�����i���0LZ��@蘭l��=��h���D�:΢��X�AaB��-i��s�i#��E^b`�Z,�(3U<u2�d�oY\�x�w)&R*`��!(\��&�Ut�����O�p�/�'��{PVe�F�;�B��nE!�P�Қ$��#�WS��I��hV��b����Hμŷ�0�\b����p
 �!����N�<����f��88J��B�����K0�Y�xx�ğd&z��Qg~	�I�p�u�%l�T�#��e�>�4����KA]�
��ӻ���3
X��r�t��) �'w�]ŗQ"(A�f�;z}y��������}2i��?z���_�I�~��Gv�s�=�b�hQ3��Ɓf��Z��ڇ�+�V����� ���Bm�q�F�a{�V�޷��};v��..�}|�Ȼd�Ν�Sg�[M>�F'F���<�*��&�S�|���U8�d�Kj-�z ���Z�#]�ڶ[7�ۏ�>�羝^:i��=e:*m� fG����63}"I�y�R��-[��V7����>D|`��SO���^���������}�"h}:&:�JF�ȲXVq�ަ� 
��T�u��$L��H��H��4b����ք��GKp�f���c{��������V�L��k��L�n�Ch��]��h��a˦�va�lvzd�B8�ќӶt���\C�<ص�k��g^�t�e���\E �IKc4v䣉|A�f��v)��r�' <�14op�:a��p��b%�����][;�>yE�rKOLݦC�9�^���4Z���<�(��pN,��Y��3�#"�;d{4h��х$�S)cq��L���)�PD+N� ���.>h�KB��fjꀾ�OG��MoCEQ��Q�!l�2��3�n*�,�3�h�2L�F��]�!8m�}��I��x�h�{�488�]�x]��nqG��-�p:Ga���|ZĊ���(nM��gyA&�XĄ��xll=@Бf��l��ٓ%-M�~UuCV�ֹ}`�����w���<�^:��Ē���n{`]`Ӻ�j��
�^�J�	�>S�������գ��~���r=����O]9������ =/ԅ�.7+G�_h��D�o%�%��zԤ�`��$}T5�)F�Z���UVI:'�V<�-�����>�����(�	�J?��DAA�Gh���2lmZg�[���9KN��n�d�X�'͐�^��Lj�<�_ȗ���M��!��q��\��Lʭ�^u��R��$������;L�|4�	oҐH�ձ&���㴶g���4��w%;>n�B�(������^{m����m�[5��S	��K'a�9�Zu�'�4��,|﷔d���(T���4j��U���'bF�H��('�@D GBƛ�a���o��z?}$\XX��X���	�p��`���h|��{����H�k��'Ew@�;]�Y87�ݳ�k��ʉ3'��'L;��~�PBk:�6�Ρ�,���y�ZW��`պ��?�\�B[�?f?�|�n���	Nj$ʒò�:4y �q(Z"�����$����� �˯�\��JL[�JL$�+Xfv֢ �0�02�@��ŢH&�(4+�8��o�V 0d��]V
B4SNG�V��l��Pf86�ժ�s���ܿa;kk���c�V����C?�,�(�v3Nٴ�DD �j�PD�������j<1��PGq�G�a!i�M�s�1�i�C�5��N��F��� ( �ϒR7���,��r���5|�H���<�!��;j��c�����}2�_���upG�4i챃��D��"�5ѠŽ�]�@���/*o�X��F��|�כV�I��G�iP \��PMya�.�<cQ���R���"h\���x�d�-K�Ck�S7-m�)�m�����"�Ȍ�3p(B{�m��f�݇�h8�Z/Z7���	p������v�n$Rv��!�v��Q�*�� w�k��`楬5�a�9��^�m�ÖE��"#|�rS���n�h�)Yσ�#�oy7^R��Q�x9������
cI��3Q`�.��7�88�1#���n�?�y>���=aaS},�����X\t�ڹ]3��mx�J9�Hן��r� ^��;�uy�x��D�P�az�i�1�[��j��+�o"���p��#�M�E��(A��)���_�k"d|��s|�ۣI>��꣰�����W�@��^O[��* 鉧�]<.l�C�uP5R<z�!��F�����S��T:�?�9�o5�&���j
���6�����/DS�a�Z!��ڀR��C?��=j�G昪"a���	�$�-�,Z�Ya�����q�q�h�:䬈�� %"u�m�,-�EGb�+M��+�H�F���q:0��}-��kW?�a�ú3�ů|��x�)K��8{�>��W�s���}�?m�'N[2��\�`i���J��E�^__���yA��ik���<�i��NU�E{��
��7Ks�%`�	I5��4U�қ��մ^	�\&g�ŢC@�v����Lm�Ő��"�� |�pY��CQ����QW��)�&A��Ng41��1����$����0�A�r1s���=מ�h�,�d�1��W�]ZG\��mF����6(ڑvJֱ��L9��2�6�0�IGmZ���4#�����M�{�C�hBF���|9��Q�灥L�9,�,�2^L9U�Q
-9��z�Z�ҹ��=ua_Ɓ蹬egla�CA'a���@��, 8WG}��5J̩�va�p�ýC�"L�q'Š����@���$�?V���Ӵ�	h	Y4m�̜YK,K9Ӌ�u��)�\3ER�(e��:��%��L�"��'Q��(.�4V���<Vc���$��_*�Ź�ͧGv�d�AC��n�IG�m���Aݴ͍��BS�k�J�)�"ģoy,��ݙC3/�	.�:]G��z�X��W�A��;_��άq���mg��ɿ	7Օ�`��|Ew=(�>(�wKa!3����S�@!>i��P�U�l��[���Y�C��w!���k=���Y�������c8��o��ƅ�0S�: ��)��0B�)]]�U9��)�m6�m�z��E��X<�������t���H�����s�~|��p��TV`//���?���!B����>q��G���=BT.���I����G��8o���]�+������������mk]�ذ1��cI���%�/D:�L�Cچ�M��a��0P�X8x+�K��s�Aj	0e+	���f�5��51@+�uh��jna�-
�����d�!�O2*U�!Q�f�l-�A3�4[O+�e�i�������^��:=3kK�s����d	{p{�������c�6{���n��Z|��l>f�z��>س����f�9�{/�>����L��:$(K)ˡ�k��,8M{��rօ�4��X(+MN�BHp��c5����-��Ҕ�a�(R��X��Ȓ���ъ5%m?L\����T�����$��?O=����$�W�z����ކ�L{�P>���,��]�wl!�H�l��oXu������ڵ.�Ek�|�����w�(�cDā��4B,�'�E\��~��K`.�lD������"Lh6n������yKϤm�S��8m��h�dK�0�T�"�)˕��g	��K��BӔ�d|C��2ӝw�4������bm�K-���L�9�pA�e��4��sk,O<m��7r\���/�����M��d��Q���N�%#xJX������*��#J�ε�wە�R�/�վ�}d���{��}vkF]���3,}�
�����L�C0ɜ,㙬%��8���n�o�ií�E�+�3��՞T��u��-YJo��ځ��Y�!���"L�"Xq)K�d6��6��^�����M��,�eҐ�ॉ�ފ�q����&qu�V4�ܱ��w,�Zo�!-m�����e��Q`�Ikl��sQ�ʣ7/�_r^��S<�fXH��s��x5pʢ@s��]��ֆvr��X�'��K�0M^��$�"�$��'�OU����\��G�RD]�5?��y�Tv�H��)�*�S�RUL��0㳟���OQԳ�ߜ�˩Լ�҆�iY�7~�5�p�{?�cu����Df����=��"āER��DBD��{Br��!�h�E8�Dc���<�Z /3�b!��!�4G<�e:i,����̴�1ųh�ƪm{���k&DsH���%f�n:"��� �E���ǵC5�A���~h+wWYa�����c������mm�1��7}v��7�n��X��zGM��  ��IDAT�i�����]�}�o��;i9�B��P���Svmy��|p"���Y�հ���
�H.cmʬ��z��%[0`�ё�4��gY���٢秭
��]k���>hX��]&��b4��a/f��.���D0?��R���ή�`u��v��A�V���YZ��� o4����͞:ow�hm�?� @��D��KE#�狣����_ڡ�:^wޅ>QBL�p��I^�G��B��������E��Ò�aE����-��Ҵ�n���L6�?�`ь��%���Q��B��Z׋嬧g��>֑�0���\<o=��[�8�T��5�y
K��#,y� 0 �C�@G��uG%���Jؠ�ؔl+%(⇷��GS�����댥��M�v���Zi��}��*�XA�O{��l���BLM���A�W�ׅf&
�0E3�R�A��,2E}�qY��Z���� �0/i�C��>�C�.|����vD{6��M���lT�X�8�,V�ǧK�Cv�׺P% ����!�������.&:�L��]��P=	��ұB�a�(nٙ9��<m1o�&�)f���8��-�$<�OW(�r���[�GY�A�Ώ��V�u�O���G���e�Io�t��Xb����Q��Cu+���ʑ�'�T^x���@���"�`i�b�CDaE_(Dw.O�8�-Dt`J�����	TD Ccw�V� �>���5�tCf\z�#|���>:R�{ָs����8����xr�Ku�X-�H���KK��!�]�i��W���O�FK|�6G��k��)Q��V'�6"��)���i�EM�����>bΡM��T�
�[J]XA���h�h�R {Î�Wjv���~��e!��NٱS�6;�������*���W�ĤI�6ϻ;�xT��+�Ui6�����|`���A�h�ZX,-��[XEW޹�&�1�L��i�	;L2�6ۇ��>C�־%�|��G�u PF�ػ���J��L*iS����:b�����вĝ�ξ�ZQĔ���#�Q�<����ݚ仆V|g��V*[�&l� j�ͬ�5��^�������Q����j�nm��Ձa��Vm����DCMp�V�"n��� �:����z�X�PRoS�\��Y��	���/$��
e1�x&uǢ�;3���SX'�����vQ��#F���hZ�?kwE��x�s׎bU�4{��� �E� h�~��keL?�_�������?���8;���6�]�|:\G{h�hGm��N���|D& 8A�RQ��T����%���p�ǝ���(]i�(q��8�4��
����{X':���	�5�b`��.\�GEWckYK-Q�鬵�k`]�+-��4l�հ�Q�b��)��K��R-(� ��b6_r�#�u�O;�ѷ8���A���0ވ��y�.��´c.��po}qK>�������]\�{���>)6�TĚ��קS�>ʅik0�I� 8+����$\������d�fS/���2曾K)�](��D��^R��$
B�:�2�-Y�E��
�I��Q=%P��������?�I��͟Bx7!�!�R��F�Lѝ��q��C������QL}|����ˇ�z���.|�w�¥��گ� V��,�0��Q�kK��W�W	#D4p)G�E�'��ĳ���P�]*��75�OT�@��*(=F+���l���"M�Nh�/ƌ���F����Iq�ƺ ���</�����_��ឝ:�h3��]4�;˶r�6�6]��tq�^x�1{���  f�
gM!��M(*u[�رN�j�F��E�5�[e���6Mͪ�P��ha������O�Ĺ��t�wՇ?��!��Ryu+��5�\�윾#�,E��OR	H�SzBu�o]�	�����f,/��Í�ݭ%m�[�ڰD�"@F������N+k+��}�����l�Y��Z���F��c�|	� P�J�[_BB��}مn��	K���_b�*#�n%9�~9���"�\L\�⧮�,���u݉���GˑN����i:�v�����)M���p���b�h�I6U�\��+[6]�>ޱn���u�,VN�o��q�Lѝ��H��(Py ��t�{�#c9��"�E�i�� �2�z�xYNt��ڤ��axO��N�Rj����A9k�$5��֯�-�]_R�b�L<�ٮZ��BH���'�$�W8+K�|Ck�����KU*���I,��٠9�ݎuH��۰�V�"�.����nN�5bC�4���ڝr;�*���B�
>�q���'A� ������w�>�����yt+Ak�D'��@���a޺�S�,>a��%;��z\��,�����NI��#}�O��X��ʻ�^�$,�XE�˓�B�A�8�o}T�%����X�1��h����䀽 ��T�pQ����e��rp?
���_�'��eV��M]�z7�f�1<���=}�Q�q�y`�N��������[�"�(D~h�`�l`^W��!����4��ОLZ��!��P���G�~|���N
+-A�E�h��_d �ˊ��!�bޭ<m
M�����i��8R`rޭó�n�#�d�K�\_۷�-����=vf�.=�8�>������-{����o�wZ���W?�9�Z:c���,~�%�@k�ET�Z��qk@�������3����6?_��<��0��.� f]�	�w���%g�����y��y� D�����z�.d��B�Mm�tĴ���]��H�pBp��j��f��|�{*��Y���O��)t�YYt4-Z�� Ƀ�~0^BƸ\�!2��tv�4���r\
+l��P��ݼr(,��|2�Z��^NRC�lh��>�+��0b�(�ae�k�A���N|
��eI�0Դ\, �P&����N�M��H`എ$����c=��\� W5���?M���i����]|�T�(!b�H]M�$s ^���X�G6:��56ji&[�:�^�e�Z��F�6 [-"+R㦾��A"C?���s9K��mTJ[��:� <��[C�O��ʋ+�j5P���iYO*�r3*���= ��za?8HH�%��x,в��ԍQ�K���x(��'ӢN�+Ey����dM��n��u�zZ���B���(:P|��%:�����P1	�`����Ҟ��X��<�����Ly(�=R�i�0��֏:�SKW���-�,t	S�	l��rt(){e��돔k��Ӽ�{��
ϡ�=*��ઋ`�Tt�+���'��(�G��1�n���2q)�hإ����x�Pfً��J��v���Y�M�#��J`�>]��ז9����עO��.�N8/��dE<�R4��Yd�����&�K��]o)��"NФ�����ޕ��8�\���I���U[]ݶ�ח���e�z�S���_��_i ��lg�b�{U�u�}��u{��f�J�U�ƌ�
~t�N�T���#_��O�[A"F���/�}�A�ٴ�b֞�tކe0a��I��y��9=���x�T�T/i��\"2)�6�?��7"��ӣ�C\m資x��i���qׄ	U��o*���L�E+�j\'ᛪ���>�2�鄬P��Ju1ЈO�$_qI��o\B�I%�B��� ����n$)H�^
�jV׺T�$7cॶ�Ѷ(`"B�-!������vP�b�5�ݑP�铏�C��]8�b�6}�NqE�G��{�Q�8�%�@�DB�\$��%N$�]Ϛ���k{�����:H�H��nG����]Ϛ�W>��]���io0	S1pMG�5�SbŘ`�������b�Q=Y$��ށt?�Z��amРh�{%���(�;D�T~�D8NK�`�<�k�a�oC,��6O�cqҤ�6�o�D��ZS�>��	��1�Q�h�Ч�B'�.�_�5Ne:�{Jw�ʔ���n`������r
���jG��L��c��!%�wG �bu���9�-P(-��T>�����#���&+�{�U�Ɨb*�;����.p��i���0@���"�#�	T>
�88~n}�r:��c*��n�����pO|Q����N�%�N�h��M�`�����$�.�2"�2���R��.�&Ir�o�@]��4�9��oUpz�wiU�A���uy�wj),;{ڒ�F4��\h�d:,��N��AZ��h�����	���A]�t*m�DT����(����	��¡<BX��?*���DRA��z�N]C ��o�+�V{����3?�U+Ο��+�v��m�ܪ�@0&�_!]��Э�}�y����m4�]���)�ݰk��֎m�?�a�0a�`��{�j2Fo�g�dQ�)����������$pT	M>j޽>j���~ 紸��' �����؉)9Rzj���1C-�-x��M�޵�'�8��Qhx��N ��=+�0�Sq+%c��|/ ������z͞S���0�r���,���Pv|�w��=�n�WH���q⍉;|W�|�Z�)�'u�z�4S���D�^OaTV1y�	F/����$�Q?��Qt�u�i�Kp.��1�ऩ��U��m�E?B(�mk�QU/���;�POOqem�
���D_Z#%�6J:^nhû������	�SG[��Z���iƗ����PS���� _�h����A�df����/��u�\�ڴ���l�,~�s�����1_'�4f�J��Y&f��˶��x/��5��8D��$|L�-�#��ȊW����]p1N�-�I�Ն*W��k���p��������#\?A�����[�px�w�+a�x���g�WL7L����|��5P��Qi���T1����J�9~��<�H="�(���(zU�WL����y^���{���0�yQ�X�,@��ʢ�9.����������.��<.�k��q��}�u�	��hNX���Ph�Aj����?Zޱw�ܳ^�f��%�֣�|
5�GYTӽGb=H���nBLG~�D�
� [����X��^��r�IkS4����UJ�3�G��R#�M���VǶ��ƭe[{�
S4;w����%[Y۴��;��-,����_�O�e{�/�E��=���!e�j���	�w�mum՚��D!pY<X�=B E����l��`����oiz�Pp�H��N�%ڔE���W�,<�P^C��������Y�q|̈���9�(�����	�DhB(@+�{˒���q���H�Lܲ:/��"@��jH��oq+c�i�k O���LLX��`U2r��{����..$4�!\]����G^0c��d@�1n�f�Kf(���HS�6���\���wpRS�i��'�R��s��%T�����'����A:�'��8V��z���Z�O�˓�
���F^w��O2�lj+�{�s�x�ʨ&�H	s.�x��4���͕zdmIH�+I3D},T�h3M^�I9*#��u	<ѡ�JOa���m��i᯵l�zk����h|X�p�q�bj���Fg���o�/)%-� rV�M�(f�b���k��Ԥ���WY�U�|Ts��G�m����<s}���XC
9T#�<����K/!:��p�'���cV��_�Cő�Gm�P��.<�;y�e�)��#��׽�Dc��P.���c�x���!UHF>�ӟ,@�`Qu�"@}���n���>�QY����ĝ��Ļ+}�����i�o�Mx��z��S?s	0�KE��&�%ĻM$$�tD�O�"��b�[�ܱ��U��¼�@Z�!�Qח~�1JsФ�^W1�Au��w#�"��,"�������������.�~�3נ������D�d4�抟��hbi�������r/��v���姧���������'_���{ʞz�	{���_�	;q�Z֛�<"���Ƨi��Çlok�:�H�-�-�1�4�F͆���#;<�X��(�#H���#6hDY[�[��i�L�o`�:!�}1c��+�6p�xۑXZ����?��cT0	%���h@���z�),pW_�&A��|)���)�l�l��Egj2�I\��V�ș8��eU;S�^��?��y��@֘�O�%lm���A�Z`��[!@Gz�4��A3���Q](�3wS�"�'���@�@�Խ�޹He��a,�曶Z��` ��i���zX���O���}�����F�F)�� '���Ǵ.K~�N�P.��H���p�0���o�!]N3!Mvܥ}��8� �u@X1�S�żǍ���,e@)�Vikj�(�����Oe,S΢ �qX2E�F�.Z �l�$\j���Y3Y<�kS/	�a�m�ݪo�������W�3_�=h�¸�ӥ6{M�Wr>g�u��M[hK$;�[o��F���#�JLե�h��{��β��;���1���>�]("猙��l���2����U�?��A�����В�ٻ�] x1H#��݅����ĢV��q!<�I����&�4�xZ�QN�N�T���w�c�ҧq{�r@tlG(��|����'�����1a��Ãl�*?��2x�|�AI��������T��p��>N��S����ɏ}�����R[=����/������ݯ��?��b�u���J!�`�K��mw�f�@3�t��|DzAԃB���J��!: [LA��0��HJK[��hA����@�U��m泙���=��&�f�Qq	6޽�B ����A|i��[Vm�mk���޼g�ʡ?q�������t)�;h���!�F{h�"��,���͵�֬9^���΀%H�0������kWlԭ�5�oS�̝*���Wd�t��F�c7w�}!\���橛6'-A�d�*h�T��%��B�*�ta�y��g}�V*e�R�`?~4��a�Rh�[0�F)D!��I�0v�s�R��SNa�lb2��f2�`t3SS�;j4�
��ju�j���`,�~Hy�s ��hC�P���dzFS���=�xGpb�ƿ��`a�b�
;�YGL�<Fc?W8�#��G�~`��joF0��{,��(� 8(���bP�y�����]B �����Z�<�-?��4�Z���:͔4�܇�G��Q����
��P|��V�/B��q�&��$¿\b��4G�U:@N�jk�LYJ9O?V"�A��.�/#���/�(.���L��v�8/
a����m��,��`x���\����M�N�vL�Ff>oi�C��"�}Uw�j݇��٨[�9�R��|�ْ52kB;:Z��vYc���4�Y��.���.Fz���Mp\�&D#�0��ѻ����!ށ&ܡOZ�]�@y��0�,b��������9�����||�=C�"W����t�0"\�JO<���׏ʣ ��<�8����λ��c���֐Gx��W���y�x��-�n�!T)����1�B�K[P�T�I�=S��;�Pr� ��Fyw����m9|/�����'��?��b�w�O��`������<	�r���ܱFm���L��a�d5 ��Qv��Z���-��Èeu{�T�
��,M[S��2������ǁ�z�{8җ8�ZN�wWmue�nݸc��n��Ҭ���OZi�m`�[�˸e�&�m�ְ��/>i�O-)g���?����6K�̩��Z����i7޿jk�oY�U��4�LAR��sDx�:��R3e+�>g׶����n�ݮì|��Y�qv�h'��[���ն�=��,�}hS0GY��� R׍�@����tn���6u~���闫-;�B�\޵R�ae��{f$��� �:t�7AI׬�h���#���}�<{�'�9{��FY8���ϳ󄠾��[��#t5�'�Y[0g1�.�Q���U����@�d)�������
�P"~t��ILŗ��]^�E\�Z��#��7n��3y9,��s~�J�ٻ��\���_�rP/@(��i��v���W�&�`�Y���igug>*�
���r?]��)�1�����ʂ�t���.i�-ntW}���F;CHHL�Q<_T8��&fL�:r|f"��`C-���i�`�f���Ez���X�0�Gq�A��]�ip/3�1����]Y���yxh�{6zذ(T
����"��KE?;�����R���
v���W��]�L�m�����P�p��^)B���ܿ��p��qO�+	;3u�?�B�L�)q�Б�>)�`̻���?+�T����.�W����wO�y��
���h�Nq�?�	��<��"�̓�<���TiCO�2룊'pJa\��%��|��(E�^�x�hk���H��ƢZL��?$!lX�}�u&����F��#�P���N<�]��n)7+�?EJ���@%�$��-��v���"��k���33<�(�hf��Ê����4��R���W/5�4b
�� �y4�;�>9��g���`j5
���$A��F��6���7����*���u�������R������ʦݾ�f��lب�Gؕ<��Φ��L�
�"M��[�ڶw?D�l��#,Z?Q�nf�R@W�ZkM5���i�:�1�/A���vl� PR��[���y݅��j`15{��������G��H��q��^B��n��tG��
��ʡ�wsQH@̶I;lW����Q�YP!Un���l�F!����Ш��nM|-���w�h���wjF.t��yOO������ +�kh��a���W湜!l�C�N�Ѿq)����XI,�Nw9uI%de�_a���n*}�
r�$X=�%."C�"X=��SZ���^+@��	��H�b�ȡp�o�.kK��Zh����tK����>�!aXq]��/�C�rt���:��g��5��7LA;I�Y�`�:UWV�C������(��Du�k�֠�Ń�>@��oT-z؁��.a&\3>��i��T��'�P��\�z�a�=�,��B���!�L)��h��t��q�����HNI�M�h���x�.с.w�r��1��̕�j�euu�I��yם���]$�'͊y��$oO����M�7���2J٘'F���:�,9𺸟�l8e�wW�T��?�=��O~���g\�>r�4Bt���&5��$���������"�G�>�y���_�PЇG.�ӿ�m����Y!B�~�F�D��k���k����ݷ��Q�Z��T:i�2vso׆��l���A�f�;���BB�\Y��@��3m��L\o~:eRZ�FU	J�v�Qe"���p�A]ꓒ��
���Ֆ@C���C����>��]��ek�l��ڔf0��c��{M;�������-�a��=�p���ߛ�u����ss�f��$���)ےlɶV� �?b�$1`��$b $8�D+�hI�)���M��7�o�<���s���:�{�J�}nݽw�V�Z��ڵk?�a�<��6��}%n���\��>���A���`Џ���b�ܽ�>��>�k�v%vn]����]�+7��ֵ�ػI���޽�E�2�m���>~�tc��iB�+�nl!�G(���;�~��ܰ�<��<ɴ��#���ۛ���m�>�;u�z���d�~�5زj��2lJ_�@8y�DGH����I�U^_�G�Ԛ, �%�hٿ�*��������Bo�����Փ�w�/]��t�_i��^�-���zL+�? f����u���ʴL�<�ee���b�,<���G�^�osh�N�����y5�y4a�ų	�����.i6������ţLWy���7o�$O~T��|gg>v��$�#��/^�:�g����!��(�'g68S�l��9��ֲ�ld|��r���(7�<t95��t����S�8����_����x�(��f3�W֣~�g���zp?9����Xܻ���<�g�Q��Zԯ���0F�����q`������{v$�q��ٟ�Ç��[�)�3��H�k�Z������ȣgϢM�����KT�ղG�t0�FN����vl,�?�-q��/��d�g|�%��P'�K\D
!�C�绐	OC�"`�E��%�<�$�s�����7n�����uf�+��S����g�7�i7o*WB����,�[�;%�c!Y~���W�/�8�|�^���`���G����^��������k_����o|&~�/��͏2�9�g��ߍ�|�S��"��E}���Uf�|	5�k�9�3L,��+��+�0Iᢆ|P�g�4�[˟�*�?�gx.Ǳ�Σx���Q>���ًk7nć>�r������w�[_�����r-v�l���Ǣ�u;���<�����8
��ㇹb����Y�|�BB��eZg�1�_?C�U-hވ	�n����i�;8����}5�f�1��"�˻����n�>
ꝣ���Q�Ѿ;X���1��[����{���p/?%�^��B@�:���1~o?��.b��x���h��!`�5��ҫ2�0]��0N�_�m�+�e�Na�w:���!��_-/ܪ�A��>�ncq����$�g}���dj�S���� Z�����W��� *�����A%m�l�2g�T��vy^M���zؚ1��Ai����P�oZ	i��ء�P��B`E��-y�<��%��u
5�Cy�*=W��x�K�E�#/I�cʘ��*v_t�����"�f�j�ˡ�a�Ќ�Μ��v���Th��7._X��#����߬B'���SarM�w��T<�6���3�~�K���,F�"�_D�x��*2���u���[1������]��M��]�� j���U�\��S�2��'����Nf��͓�2��ls�a^!X�>/e3�y.�ɻJ�C�2ެ~�'M3�N�� ��}"W���r���f˩9����,ܑ.oJ��Cx4Օ���NUvjL�u��`�T.K�����d��4�Ә#�x�x���"��=4�Sr?<EL`���I��Rw�c,��|���I�uU).w����r���\,��w��/�'�0��aq�7*��n#^�����^�#��XEkw����������K���c��u��e�ޏY�(Z0v}Z�����?.�������8�md����+�,�����A0q՘����[���w��/��h���wb6x�x�(�[;���k�޽�x�k�ç�j\�݊��w�b8�������moA���M|��oţ��tT�\�FyV�F���s��fw3|k����j�C�FNם�A����,�����o2��}s3�6���n+>����o��{=���yp[t���������T<�Zz�v�������7)x猺(;z�(��8�Y��
��KfJOGF�t�>�����y�%����w^ ����9]�E���h,�Q�x<k;<�zL��:�?��{O�:�E۾U����z�/\�@y��yxO�@�;���?�깆�*���蛃c�fH`�T>Ypzt�&?x�rU�e	��ro���t͗l�����^#-i@��/�Q����^Ӆ ����Z��.ʕ1�})k�J�r�~s�)��>�4t���2�|*$����񗌭�����T��p�9iHg���j]�Z���Tdc�C��x���z�M�u��+n]����K�O�1Đ��?����+=���F+Z{X�77b����&�u�1c=��j�$�&v�i�S�mqzWY�;i�=~���I"c�H�e_�T��ϳ�ȹ�nY���F�[��~Z�e]�%ad#��sٸ�ԛP�����γmG���S~��_��h��WY9���dN��r �$�o^�8�w�U�?,�r�L�g���`�s����|.��D#������P�dQ��C�B�g>ԡ�T��<擢j�K"*x�~�����g��\ɭ@��hӸElq��W�1����7��?��ߌ�[_����)��K���f\�m�F��YP��a.� ������R���ee�	5S�L�'�0М�![b���7�������Ø����5�叽�����՛)@��F���A��/��t�ݍ����8�����s �𪜸��E?�~�=��n3��P?�r�СR��oe:B2�����^;z�F��:������x|x��o��H�t ��=
X�"\x>I&��dDdaX�d�����`O��vt��)M~R����d4S,l^ʬ��˚J�<ʠ�lE�K��`g0V�eq��V���f7��ݑٯֱ��x~û0��(�Xӽi%z�D��h>�����i�J�M|���-�o�m8�����<����oR�9�F��D��A�Y�*��<k��*��#�|��<�jNI#�&�G�6(gj\��N�6061�>v�j|��v`jDO�6�G�3&/��gC��5B�� }��w��>��υK��׵<� �9W�xX�Zt.�؃�+�7'n,�1��T�[�p�o�|�e��ך[�p��v)u����}�[�'�C���saύ����L�x�����E�����iT�g�لj���ѼB��B�lƤފ!�\*t�W�����!��k�����,��4�)G��|����E�Ai��� ��ϴr+p��k��ט����:RId=�$��yI� %#��QeTF�Ǫ�JD9��]�'���S� 鞹��>=b�K�Y¼�H���w-�3��sʔ��v�O��sK�N/��4����"�H%-[�����4B�����<�!��X��$��3f�@�LL	g~�t�����h,j�-vi�����0����[�ۿ���{�3�k�M�������TɼZ+�h�
g�v����
��Ky�ܢG��.�T�L�qx|���{��������[7c��GZ�g'�8ƣ89e �2	���z��:���Ay�[����wmt��"�⍷߉��F~[��r#�j�P�C4�pԏ��E�j��p
B}9կPN�b1�	�f;�������rԵ6��i��+˘��W�e�tr��^�A��e���p���Rh.�Si�jJ)�ԖCR&�J��#�ݙ���f���23��l[�,�}6�h�<�Xˍ�x`�ַQ<۝�wP�2�p�`&��y�Oѥ����*}�G]GY��j�3�f9��r��{��_��\�<� 0�obU�2�G+�lЅ3u�|�`�ghZp�!���U��t48�ò�V<Zk�.��p��|\�ӟ��}�
+ǓD9;T�oRA�|	8��O���2�ay�,�4���g{�w�(�kqk�?���C�����0Vj	/8�C��ӓ)�����z(܊�cC��^lY7|�!v�BhN�|�E~�����m���Q���%��P~�w~���9��#����'���z-�W֣�����L1f/�ԫ�_
u�kH���̦`�*^���|g����7�����p|؇)@	�ų;���Vz;� �ez��'jt�	��/I���Bs,Js��X�K<�L& �"�޳��Ø���IykY��K�\��S�<�T�6����m�bl�T*$��&�'KʓY�����\Z�����E^��2�����~��Gm�e?Z05��\��rc9����SS��| ��kU�������7���o��wވ��1��<:���V_ϥ�i)��+�\8���C�4��F-~�M�ݎXG�������'q����h����Y\�<�Se����[{xb[x*��:��9qg���up�K��8���f���Qi5��8�<�O)�~byR�-�m��.�֓�9TeӬ�	��^���r��;��d^�:.X��/|K[[FB8�UNtIާ�O,����?dIA��T͗���R:Cv6�벙��j��-��ʆ�y�7�U5(S�)$�I��}�����2,3���E�h\�T���h� SEU�p�T���R�%�"H��,y��H/0�#��"M\��h�r�j/E�B��(�]��u�-+�k�iyuI�Oj8଎ �J�����ݹ��b<� ��e�<����:�m>�����
Ȝʳ�@�A�i^�y1�P�<�xn�����O�� w���`>�P�R�<�
2y���e=�	*�^��L"_ֿLW91vk����F�mal\�FmE�j�ٯ�LR����<k�~2}���(�+'>���*������\h�$�Ol
�RЂ)پ�����)�P��"3\���B(���)����Y+�OJ��k�kL�o%��Q�bY�P�K��e�	��2M��I�#���8�[tun�L�������?wmX��U�T����2�
TCƕtIg=9���e{'%o�����<�
�rL�i���/���ǒ���,�g9D*\����JN�y���IS�/G�h�.i���$~�7�?�;_������6��Et:�����O�Ŷ�a��I��PpJ����&�yH��K�����#ೈ>
�ޣ�q��}�$�v�b��gq���?=����ؾ~5_:�X��܈F{=�����	�D�jM��.x��������ލ\�):��[��I�d��V����n���u�O��xV.p�{�?D��b؏iC�_N�&�	�V�iͻ����<�\�ҷ)\r H:��WJ���avq�t~Bf9A�
���w�����_Ц-ˤ%͑��r�!�<��4kt��u��n����8��#���a<~�aL�c��X�Q�x~*��N�����͏6��/O��I+�mq�k�In�;�KeS��c�~ۛ�V��(��bKq����G M�ۥ�G�<�?���W�*,��)��+��_^&�(��F��3|�W��/Y4R)�Ro �1?�H���%��ȒÖ0Yo^%�P6�&q�R��en�/m�2^r)�U|ڽNL�s̪�z�<�%Jg�O��Ԩ�.��F4v�Q�8Yl�b��3»��3�%m�J�"k��e������|���n�eQ��dh�R)?h!���ϳ@J��Vm_1V�!�{I��.=E��J��Gy��,WJ���y,��0�}�
�}o�V2�Q�A0�\�`W,��}���7��K���SBXn�r�Y�Ўe�U^s$M�!#��QR-�qy��P�N��RF (���������hy��So�E�&5��`�����y���~#�����8����4_����B��ã ��Ah*/� C <�*�b,WsǄ;�?���c|�4>���k��x4�~�`ⳓC��Qtwz�Nx��۱�w5N�O���;���o��u�+Ҏ��Pf��w��ʴJ��K�����Y� �:�y�)|�M,�N���fz>�n+������A����>֠|h F�{t�4�˷�����\4�+�I$�!�-�iu���B�.��_e���f&��j%Ua��S�2%x��*�ΒI8�ͺ�Rz�>o�#sp)�v{͸yk3�].�#|G�i��_����qx�$�[aY�+���ʪ���'K�IO��,[�/F�R2<�Mb-WZ��i2�O��V��}�rϗږ�+�n|M��'����c�>�ٝ�W_�u���S���Dzж�Р-f�=�7K$C���+��Kхi=�-JZ��A�s���ɀ�#�¯��Җ�g�����n|�~?.��P�p@*Oq�����X���>�-���9���u-��W!n�:-oZ��k�����6��+��_ي�N;��[w����L����0*�@h�'%4NZW;Q����͘�.tsz:�)BiӉ��9��c��?�����\�ezs47_ ^����F�t�#���_ǉ��_ �g�����{�Y�Dp� ����i� $�2�̟xQ�_��`�3�$� ��=
�Q�R�:=�-IB�ɯ@�^�9�ˑ9��c5VL)p����A�r�W+]Vp�3�˕+׫ڤ�2���"�s̖ˤ�?�e���?�i��=��~�+�����ٽ`�8@\FwA��������<\P���Z�~�\��E���bԈç�����/�~<�qB���Y��:(K@����={X�~�$�Z��2�.�O�~���o|3n�����ػ��e݂
P�Χ���f�/��b*����f죸���Ty�ƻwƣ�1Oc�{W����N�-Ӗ��v�
ׄ^O��L�hcc��e����m�U3����2��w���Wc��8��bq����-a�lvb��zP`Gw��8�A��^'� ���y�<����I���9��zU<W�ɬ.�M��2��y&��2�J�̭���s.�����N58X����_�/�z+��x��I�Q�+�.p'�]ԡV9|"9h�NM���jP$6ĕ6; @򿝘<-Cp��m��^m3x)�/����\���p"\"���<G�ٳ<į��3O�ؕʣ�@ �NX ��8��gue���ܪ���w0�mʯ�	n��ۅ[�%�
e����g������֣/��
ʣ�e\���G�8�Pk�]��^2_���u`�����c��u��m~Yw ���|�Jz}���Z\��{����C]{�X��x�q�k<B����i,\D����l�����y}3�[1�����0�)�+w�(\��� �<��Ӽ_F���>d��F�[~T���<�_���ީ½(���|�l��WxX'Ǫ.R��<,��m.�1䏱),�8'���(W��,	VS��m�>%zI��V"��.�H�	+#��b��{�r9_�*xd>�Y�J��Ea;����\����0L��BJ�)�����w��S|p�Ő��+W���a��Kn���!N�%���t|�i���<����;��55�+�J|�J+^{y'��уx���h�`B�BG�ܱo��z{?֞�|�:��j|����?��>?�ß��hgg��Y�=���V���ӂT�r�=�t����$�=9�?��?�?��׷6��|-��_�g9�T>�=���nQV��0�(���8?:�㣳-��A���Y�=|�ylmn�g?(�ݸ���Y��_)����}o��'�g��n6𸶶�sza���� 8L����88����������ߣrR�n���zT� w�/1(_�ĭ8�ފwΆ18���ݣh<8�+�Tx ��)�m��z�p�}�n��>D:^�)^ǹ�zx��9�,����\%.���S�K�d��9B��٨ru!���ޅ�*tFs3v�_��+��E�;qa���k?fGѩ@��EL 2����	q�+�3�zW��s���a�-}����ܞ�~uS�z��s��5\��GZ���P.M6g��Pf�<��,��3�L�I�3���xT1q�6�Da��'ޖ�i��Bdp =��UzX�2)�E�Ё���0*yҰ��|�T�~�������1�(8�kk�G���
83� �L�\5"��m����]����z�]�})R.���񬜜\�����?�W/�g�ky�..@I�}�g��f'���x�˯Vğ��8�/2�a<�%��B�,�A��;�kG��\���'���S�dDF�c��[BB3�W���:�TT��%��s
-S�P��g�x�#� o��E��2S��)���aWXw.o6�ϫcE��#\�]V��[zYJ:ڮ�&�g;&!g�q�s[(h����פ����l���!;.��ˬ�bΊ!/�G�%������h-	��%Z���g�����{������n�"� �~M׻������A�����P��pZ	�}���wP����/���C��W�U���h��4����+ƒ����,^'	�π� ~��������#����r�ć>�����!�.��\=�W���!G(���s��I����"�(����xzt�?ޏ��}קW�]��ׯ�6xv{���D9���h�ҹ-�^᷹������(���flo��ɸ�C'�(��x�;ZG���y�w_�63�ns'&�V4�K�kv��v�Q2�c<�وA<�.��RV���cp���g���禤*���$�v,̐����F��]���I+M��xɤ��VZSNfW@��L���i.P`8zd:��ZmDe|�J'��Ɲ�Q�qr<�ٝ���P�(�Z��i��GdNqX��>�N�p��֬��2�~�����e����ύ7	��ڀ��^㾦�����V6Վi�<���m�������m>p�G�-u�e{q1�K�4��m�e�7D72�s*}Ap�=���^E��Z�)�Ϧ�0b���zǍU��9P��F�@ƌj*���������Zt,�(�A��4�!��gx{�����q]B�w���#]o.�O�F���l����e*�:u6��6�ze#&���0�s����\��@���<Qzr�+F1!ӑvz�1�
F,y\�!ߎ}�	 eLYj��\*^��uw
��`^�z�.'y
��x@O�$�rV�P]�\f�V�T6��3�O��	�U&i�� GeI���M"�s*���[+�o�Z�HD�3"���1�Z�a[� ��g�X\���8���O����v2@��� n�g7m7��ȗ���Ac�	&��𥷴�T�g�!�<�5����<�0��;�<SD���v�Fw�f47o�ӳ����4���(����FC��(�/�(��x����ӯ+�}��AA|����[�p�hC�~D�L�?�ӳ~��<|�O����4�_}���x��ø�� �|=��K�߈�o]�mɆ
����01�Xv�te��A�nntcK���Fܸ�����;CxJU��"Q������B0�CHTCh�`�#����.@��|g���K�%B��<H[��ZMN������!��-.9n#[W7"v�c����'�Q�.�\�`}�c�f�K����V�ԛ�N�D����9Js��@I����%��5k�48rn\ށ�VBC�F�O��~`���"1>=��*�S�A���l��+����Ҍ�s���H���j���.�L���0�%��V�Ҋ��`�䆏���z��1���S��WB���y�δ��s�C�)}��2����G�/ƒz,�K�'B£��ӹ�e���h.+��b��N��s�?�p�H�[X�k��֧��*J���^�x`���T���D|�P�`�ez#��=�uΨ��*;���-x�Qŀ��	G�xt��x����t71Ԯ��q}+�?E�/|� �e��p���5t�^���"+�)y�����_el��oP����{��gt��D/�l���X�$>g���{y�N�k��K�^�>&�E��/�N���Pz�oR� W�����d�
��
��;�s�q���O��g��4������ ��ѹ�D�'���9)YNy)���@�M�R��Z��O�=9������Չ��UH�j����[pp?{6U ?�(?���Pi�|��w��/���O��>5Sb{-~�j7^|n+�s�N���iZծ4��LS�ӗ��Y����o]�����D�_�͟�+���0;Xa�����	L���I��1�ǣ{ocT^ⵃ|jg����D/������Fw����l�㧫U�N(̍󋢾d����p�c6�!�Q��i(�.
GoL���\����q��?:8���%���Iútw��UH.���j��5�X4p���{w�F�ƻO����oQy�46n���X�뱻׉w������J�I��L��G��Ӝ�jbq��s��M�|p�β3�v'�*�Wus=�i3f��ӧ(��~4�`@��)��5
AbieǗ)��	�BV撞*�|�$���黭�F���������x>�ϧq��"f�ޏ���� \&�������]���r�����K��::�'v�$��G�Я�g`��~:[�޲��$�	�UЮ*$���9����H��E.M�TJ\�6W^*�\R�ȡD�-7�HU9�d����)�[v�?��gT\$H�)+�(+]�ϟ4ϊ�ÓB�<�t�re7��clN��|�
]0)́�?�RH�a��K�N����7��_.�W����S�'���e<4`����|�z��ӨO�9�U�lF��V40�ƽ�al��m�2@��{�0��%��L��8D���%î��^&��%M��IɃ\@��u�������L��e�t��(tF��&Ƒ5�7:�ٱ�x���#�p��	�Wɟ塃x�rIX/t'��N��b��>���F���:ҥ��"�W֛?��g��_�aƗCŰ�3�<˛<9=�����;_�ȼܛ=����F�xQo�?��]��V�cxpH{��?�y6��F�)���ow�����@����G�/��ߏ�?�G�醭����V�t{'޸�~�y�1:��Ո1h��4��уX;Be�rYc'~�����;�g�ʞ���T��p�]�d@^��ܿ�F�?~0w����18���ųx���ccs3��p��,��oi}-u����
`�+i��S�B�Vǝ
j�Ή�FB8U���3��`��q�
i�75��� ��NԦ�Ϧz(���1䔅�@�`���x���q��(������?�ŷߏ����Vl7��w��V3��{�щ��'x2�8�wݻ�(��h��#*�?��,d;��s<������k�mFm��@���c���bqt�ӆk(�����r%�&���2��"f�o �B�K��G�٭Ň_��Wz���8�_L�~�� 6`�|�� R�i�)k�^���s��I;݁��p����B��	Sv�)��p�;2u�� ?}^�y�Ni�Ih��+-A~�iQ���mŦ��׭�N�@�������B^�n������H6�e]PF�]�D#h��$Ĕ?i+
S�W1���;���h3���joѵ	/��\ܻ� e.�������X�4�n��-�_�+�cB�#)J��6A\���F�[��������{�n���F��q�sm7.1��(��m�����rI�"mR�s��Z+�f�'�jz$.�b��0On4��h�euB�L&r�ǣ�s�8���vȗ}u������9�u��"�s$|������՘L\-c�(Z��L�zE&A�|v�L6�%�1F��v�^�ȩRq$�pS֤R��>�gE�G�"�^��eR|�i_!�)%�J��6P��9�K]�)ͪ�|���OtT�����]�X�#!m���o�M�2�[�W�蘭��罣A���D����b͈����n����1���,U��	��a���9�+�n����K�}9�ֱ`).�eY�3(qE��^�u�W��r�`r��Zy��;<<��O���x��$�=���'O����q���ߠ�su�%�Dw�X��UK�Q�8��w]P�ss1�9I[p=E�-�DRH��>?a�7��R_8u���Y�����Ջ��8:<�wĽ���I#4�����>��j�&,+�:�]���1h4sW�1���j7Ay����;���N�1�	ىp���t�P!��ip��!�o!�L��� �#���T`�\��IG�me����"����Z�q�'r6���mq0�y݉��+�_v2p<[ںU �A9e�xH�	���Y��ti��9���s��8��c�������m�B�7��_�:φ!��k�zo"����u�����i��kWbb���|j�9}r�gHX�aџb�sM�>�X �Y�a�"�Y�_�@pqF��gƙ�p�Np�s����VUsiH]��Q��s�����-r�^e	7�Yx��������=x�p�#q3�I��_΄��֧��L�[O��$XCq�n �i/��R������a�"1u�=P���)��58��v���� �AK���=�~v���
}�0�I�]�6�
m7�jc1#�ƌ��P�;��O�B�M9=��%�Ĺ�i=K��R�B�^C'S-����4�my��	7a����g|*���3GQ8૑�ם��d��|yp*X}p�p^�����q��"��7
�]O,�e���A|��q���hH�"+�F-�|T���w�lF9jU��i����N'��Aa5K�V�s�f\�]�c����Eji�W9�J�"��E8dc����]�����c��p�Vn�ʵ;�����1�8KkC/d6ᥡ�G���n��H�Ѣ�jE����R��[���d�{͵���6�0�L�0
�KʌP0>K�%�}�]�WO��Aٹ@�2�Ġ?����ci�6 ���y��Y�C��Y���Qt�x��(�<:�(�;w��{��w�ޏ�'���oܼ�G��?=¢��f,\����n�����՛q�Hq���l�SЙ5�O.�L����2�f�3+7�¹2��/�(!�\w�uZk�p�`Y��Q9�+�d���:2N�
K?kQ��\peZ�ױtg�#�=�!���D��j�7���eZ�MxɃ�-���E��nFuo=���|(ߧ����{��x0���I�-�����g��dҊ��2�A���A�A�n�q��v=�ŷ�s� ��	�p|xg�#1�"��!���íj2�6�9�-�6������V�:�Y���G�)�������� s�JϾu)�B1ar^8�Pำ��]y"Eʃ��A�T\�=�s��ŝ8%�¨3��7̸!q�)G���ʺlw��<
���kF�>��������>+��.�+X�+#p ���:������r/��+Gɑ���ެ����(c͛��F<���Y�~}-n���� >��zA�u+;�K�	���K��E0���S��E���F�J��b�8�0��N��e	9&�6k3���"?{�έP>�:�|����ի���<Ģ��ؖ��dۑ�s�Y�@�{�����$4)�m�y�fy'��)�XJ��f���y~RC�x�j������P<�?3NϹ��w�?�_��n���}�f%~�j7>�ʍ���o�[X�_유��z>�w��>���%�7?�7�\<������r�����?�7���`�Ǖݭ�z��y�ʱhq�?z'�G��s��Vn��f�Up����]z)Ʃ�!Jc��0M׀�D���_�2�8ϩ��X�T"(�}_I/�gJ�ӣ��;�\�� V�N����@Lg�|z?�i�v�:5��
��n-^��+�u������x��;Ȉ��w�U�;�Z��l�K����,���Q��;�ޝ��j�@ʩ)_��sZ��e�����\F�`�6ڬ�n9���+?<A�>����E@����-�ѓ@��g�E*�6�9'"H�:��}������8��Ә�q��n]�+��ŷ�K�2d&!����{ށW{1���W��1�y��A���t$x�����cLLi_Z�'�%�7G�"J:Gr������+�(VGY:>|��3Ct���}�zAg�aj�H���G��B�tY?�+9�i
��ӶCg��J���F����%<��%�^��9nҪO���0�7��'z
W��f���{�B�*�|������A�����푼 . (nD���j�F�1 �����uc
�k��ߴJ��~M���x���Ռ=���>T�R��� �4���p[��d��e�L'-��e�d�~zk?�����A���|/���^�5P��W�?���&}ݦ^���=�7��Sq*�o�)�4Ŧ1X�(³̈́��
�%�\�p�'�(�.�_�Qۼ���U�5���O�;(�3�v[?��%I���Ļ�5�wWy�������Ӳ�y?(�p���
:���#k��G'�[�����?�������ϕ�7s�ߜzK&�����f'}��]��o��3�?�ï=�2��_�ދ�|=���y��c��8�������oq�����`�>i������+_�/��O� �� �ܹ_����[���蟝���V�7wb�"9::A~�������5����Kk
�L�ڔ�uzԇ׹=�:����q���v���7������0�]8/	����6w1��t:���#�O��K��� ��Àw^��2}=HxΠ=�	B��^/n_ߋ��n\ݪ�G_}>W�w������dq-~��'tX+6כqc�Ͻz+�7|n2���S���*:ȥ��|�-M��3�C.(�p>ե���qIp�
h{ϖ>-bp>��ӳ�����)HK��w<�̜R�0�gG�̙r3�O�S��>r#&{�x����p�7c����=}ӿ��%Ë��S ���}�ۡj[���c�9�����i��?���y�`!�-��m�Q��M�2��B��/��P�e;TDE@�S��D��se��gx*0�PS��1��\�в�
���� #]ϥX�ū����hY0�Sȟ���g����W�����tu��V������>o�F�
]¾*�m_��_�EL�$J�
x���-U��OO��x��3�������������<�ݫ-��V��bbt-�$2���ɛIt�Y�#*5�0Qb9�����Lg�[�c%<=
��%�-L��^h&�4D�w����������v%������'��w>?�ٓ�n?��1n��FL1B|���=3Ф%��(h彬e�q�E��&z�� ^e��$,_�0~��6>�˃�Fc�{�9� �r�ޗ�_��y;&���ư���R���4���}�{�{��-�5�Kt�~ ���>�]�F��	��W��b�|�Y��A��h��*�x瞃��HFE���gю��NQ>��7ǿ�w���xR���#����W��ｃ�y�w�0΄�g`U��� m�0��������+��/�'��������8==��ē'�q��\�b|��uqVS�� ���XkkM���*�%���"u��1�`V���v�8ToĀ���v4�(�6<?��b�� w�YzHnR��Ho�%��<%W����Z��q������p���m�Z\A���^ܸ�W�#�7;1�T�͇���G��݌78�X���F�xe;�_�g(�7χ���9Fy�|vT>��tln�B?�����a����&C�ؤh����uq<����\���<ڮ��]~2�e�a<���R����������z̮��]�'t2B����ͣآKz(��=J���`��+�6{��r%�ьc�d=L��3�{�?��Ƕn9|�65?5�D���>�./G:��t=VAr) �;e�Q$�R���� /g��u��Z��%}����I��֞m�>~��> �2>H.m/�E�Y��"
5�������~����buыa2���z�O\��8��\mG߀�5�K��⊺��I�=Ǌ�zQ3?�)��0�7Q��(�c3w̠	�\���7U�@7FC�.���\�T�,D�tP1�T��/EE��ɝ��v�A��&/s哴]Ex�P$�]���3(<�\CȻXg�Cl:���1c ����0��Ň^�s1�z=.[7������hz�������
u�S9�q\f�R��"�f#�kn%n>X����tZ�v���Z|#��1�}>jW~,��[q
>c�O��b`jHq�jq��������� ^�MW^r-ٲVcz��
{Y�d�dg�^ 6�5_� �n%J*�[�;dl�=�a�|ɔ���k�}�������I��j����d��o��0����i~��ٍz����ya7�s罸��gS�iZ��S�?9�řb_F����F����������؇�+,�tF����k�OA�e(I�ym�*,���`"�t�!�Q�l�g|}n���ڵ�Qio�pr��ݍ�C'ˁ#ٳs����Ӓ0��+�w�e�|Ι�{/d���~ѯ�ۍ�F'���X P��i�b�{���͘M����z��3y�e<���x����q��߽s�ZX�d:���FMt�̐��[a	̢w����N�hu���^7�aO�3����qL���L���n�_�_�4Ӑt��q���zK\�r�>��7c��w��x�w�c��il�S�+ޔ��"�e�܉����|���~�3�V�$�����O�ѿ��~p]x��ת�|j�\�-;nb��Z��1��:?8��~$ޮ�9)(�cN���9m5��-�R�lKX�M�f�e���>Hz:֓��s�+�(T�40{
�bȘ�4�$AA�p�/�'����y�̓���F��uǌ�4Q�m\�nۚ����A�Q�|z{) M��ußm=U�ȭ�������?����M"k��W�/^)�m�g���AeD�(˒�dW���/*Y�6��/gX1���"/l3:3R��J@�AwSY���v��OQF��������1<�N��_�����*���8��ogY�.�q�À��9T)-�Q�Nn��v�
��^m2���3å�<�"=`���땋h�ߎn�'�b�~c�31��E����G[��]u-|?F|��ؚ֬�P�(�A�*}k�4�<Vg�ե�2�dI��G��M�k����QA)���9k��1�?L��xԈ�����\* ݐo�����.8�կ�}0���S,�s���v�{V�u��2����Fq�i�o��|<D`�U� �AQ��������`g�kq~�k?h���1�R�M=���lp˅��nޏ�o�ڂYɷ�%l|�x}�O+&Pa������+(�-�S�����,rU�``�U�mn���[3.u6����uB���7Z�S/�/�v��Sބ�B�!=ҟTb��u�	z����ݮ���v�3�O\�0����)^	����fZǹ���pIK�Φ`K�MR�e�D�v,o�s�ƙ^���v�v���X3~�Z�R8%W+�`*�)ڑ
@֣��y���vvP��F�M%��b�x*m���sT�X�8���#8���:��*��<�#<�s�泣����*���6��hb�T�:X��;<��WyV�T4�zl�����숰%e�!��C!"�NaY��z��xKXy�{R>��Q��U�p�[QI����w���g;
����k�I�Of����g�	�H���q�=/xVЛ��o��SM��{��!,���t�Ug�����*�,����%y��AZx�s>�Q .a�6���^�V����Uښ�����K��T\�1aAˉ�E3�!Zo�徾J0��3Lb�t1�6w-���%����<��hҋ>
�ok��ּʾLV��'v���40[�w�.yKF���h�?�9�HFc}^i�p�����vc� �NU9͜�U�b�q��� =2�<DZZd(Y���ϔ��T:��-��eZ�/7�A��{d�E��F�.8���o	�Z;��@�yF^Wz�e��{����>��/)���ϯ7rc�㋳�N�Am�oZ~�u�6QP��0fV�`V8`ɺ�-
������m�{���(�1ɀ`��|r9��$V�=�:�[�-,k>���H�Ӎ��n4�w��]�%���5�����N4{�h�zQ�z�¢�s3GB `��-I���]]o�ֹH��I�J�Բv����m{)]� y\i�lף���\�i}Ô3F��k.u}*�h�[&)I�?t��I��HҖ<�̩�}���9��8�+�N�+H����S��B�R�U)X�Z�� ����n*�K��_$<>��������J^y4'-i�&k(���A��q���?���a�Ч�f-wOolv���k띘@o7M�+�*����Fd=e�����[葏3�A�i^���a\�j�+��+��)<�M>����	k���u��N:*%_�Ϻ��:k��������/�6��)��^Ez(���|�}��*i�+A���ĕ��!iBZ�gY>{�t8�����<��r	���ݨU>�?@!�Ax�z��T�����9�S��'���R0�2�
����ڲK����2��8Z�����Z�!����R#u�Ӎ��g�LC���|��L�xA�9�q\�q��o"�-�sIwc�Nb�O~�@D4��2;i�&�m(�=�N�#z�q�TG����Q�+�	9ޕ��+��2�+q(��'x���w�����xV��\&e�l(Qr�O∓�O���U�dIK��6���4Bfv�����_��;G���o?��>6�������J�j����e�ʧ� ���E�B���g6uH`��S?)��>�Z�w��@ho<#�M�u@�8�^oG���.ʯ�ν�׺��.�(�R!�����^5����zl���8E(3��8���^C+ڝ�]���*��©rv0_v\Óq��5���]�3�{���>r7a��5y*(�z�"�Eu�]����%�0E��RסǤ�L�!�����Nt+#�����Y\���-�;�e��إs�NQW:��%�� P���.�N^L1&��t�@0@8���M���R�Q�}ƶA��h�)����c?$���д�9�_r��V�3�� T�t��V/�b1��18�{ztճ���F�7�ѻ�����SC��Cyߗ�O�����{_�L���E��ȌWXg>q"�њ�?�a"J�\��0�e9�0�䄕��|����$�^��]���/e��Ȱ,gi��q�g��w9�\��u ���l	^ρ]�S^�x{�4ېJŸ�O;����[i"^��?�J��~��_*4��Y�\��fX�˲%-���~'>0G��E(gTJ(�2���ܤ�i� ���+d^�fU�y�e�����\8��;X\҆�ϙg��77.��y;���̚����Rȋ��&�+|k�
HE���i�Y�xӋ���9/���Μ.�Sx>Ӛ+�/�/#J;����L�u˗ڒȉ+#S��F1����JF�7'y�zvm���U�,�M)IUKz�K�	�|�-�`��C-ɢ�ɮ[�3҃�,��{ϱ<_��7����_��o>��z��[��K{q���x��Q�V���įz.����~��Il��,�{jv@�`��l�M&Q #�lpZ(^��ì
Y2�8��_��.dpq�>�6¼����ĕe`�O湀aqя�h���L���
�TP�B�?�Lѝ���E^][:��}���H�C�;�F����G���G�o�ϡ�ٌ���Q�y5NP}J�����qԞ�F{@^�AN��|��(�o�89��!]n��n�=R�{~N��UW�B��g�Ø<8�͋il�e�iJ���s��FdJ���7Sz��x��+1����8\ƣ�gq��Q����s=d�l �	�]���-����6�����60�_�	��Z�gq�s���^':/\�>k����M��`)��F����\g륏������7���.IyX��Om+i���r�!�Z'<h��O�N �x8'x�[��]^��]����.ә߇���/1޼��%����⑃����5�,�)*~^f�2�VB�#˓Tn�݌%���@�ڲ6K�[��:�w����x��e�7�:4GOQ�4�I�UZy�b1*(��b�D ǭ�\��$����Sm\�3Vf��%���t���JF�����g)�Iw�e���˕������W�^�ͦ��O>��-�M�!��F=�r)c.��q�߃���I�$�OK{j@a�W1��-��|�ۤ9�D��Kӥ�3�Q�&���a��<l_�W^/����{�L@�e��+��;�S�,�#�WYp଴|��.,��H�K��ݲ
��u�h�����_�{߈�o>�PS�*�F���v��w��j�,��n�ۈ����R��A�4����%"WP١�p]��80�ˎ&����HB!'-o�K�z��UG@��:���pWpʠ5�x;����T�%~���ב�8k� ���ގ$2ӊ>v����yZum΁&62��\�,L�ԙK�(�;]?>��x5A/�֪�ڵ���v;0祓�O�#��Q�( :���%��g�NFI�b�<���]��*��[���M�����2Q>��~2�]p������d7XG��<*���~���1�����t'q��<{�8���.mO��-���d ��w�:�­���t%ރ&�M��x�=ھ�C��c�W��y���]��z�JZ��δ?�S�1�a��gs9�,��0�P>���5p Z�m�0���s%��B{���1�\]%���m�Ϝ6����֣�� ��H������R�RG~���ړ��L侴'�͐m&��P�#���M(m��7�?�y�l�c�Vym��'id=K%���U�R#�c�(N
~�&}8[�!�7�U�0q�!!�qΚ���|���f=�����L>�_���9]�I2�wj<�����ί���b�����%`՚k�߇�kȑ%�$5!��:�X'xK�T0��]�ｴH��F�?�b|���|�Q����[h���k��8G�(��.R�q�F�?��Ƕ8F�k�(�ˣԒ�V��{�%^��˳�rdS����*EX	�����|g��9!��`��c:Y��Qq�sf|�
]��F�Aļ�w-c �ȎAq�x�k�;��l8DX� ]�z�ׯ���;]:����3i��M/���hz���n�l�ջY&ȷ��!{�<�/�ֈ��:Qow��mE���4��>f�}#�e�c:p��^U�Q%?Gc1�/��W�	�n���*0+-�(����b�53R�YkDNlT��5�_�������6�m��۬��nZ�X�L9�u�1�|At��Z�����z\�h>؝�/cr1�>����,�t\����Ѽ��RڌI�cF�t��|C�� ����*���@�y9d��H_�}l}˲ɨ�ja����*�Y`%d�@���Cs]|�J��H�Z���V��=��/���K`ͧ��K�2yQE�a��́�ӈ�߱�2��B%4�L�����ܕ}�qʝ
F)�-o�m[7�j0�&
��26����7:uT@�r4'�u�Q�3W21���g��2T�9�Q�\�r�L|���5����(./��� E(�ޘ�����A<��t�L�m�k������(����'�m�]�U�yW��}W���0LQ�
��V�e[(Cy_�L�и�P5����)����9[~�TRXgM���ԙ
�Lup�0�s�0��o#��b��� 1�b�������C��],�B3�E����K\���`p�H�O�Ҳ_��И�.��b��D�mS�s-�Xڢ"��������Rz'K�f��/a�xq�*T�#�/�:�V�i,i��Q����&�N-`-�#����!^g)ڐ�a��rC�|v%��'��e�lŲL�y�iY׳3I#�*yJ���?iZ���Gf�����b�d�Y���\!%ώ9�7!ms��G�4���p�H�$��l%�C�u9�4�<�A��� "���&�NUޖ�'�r��K4�$��'��x�� �rܸ5�i�\'4<�5t\��6"�K�u��)gX#n��1C���s8���e�)֗eȫ[�3���A)��'��|뮢H�v6c���O00l�6||����M�t�x(�k��tkz�C�V�}��9=4��{δ1�G����ħ'�^O�Y��Q��,�쩥ȾO:ː��8�s�����b�̝A��R���]²,���^�����>���1��n�rJ��fAr����.��Ms=�͗�dL��*(���a�<����7��Ja��:��q*&���V�Q&�
`�g(�ތ8���-��{�S3&�h0��`H�;q G�QT��*Gۗ�S̢��Y����76z��[BO�5����<?'��R��a�q�a��}CC*g�EEY��Wcl�B��.�O%���+Z�o��K5���RتW��
a�VT�����.i7Ÿ�'�iu�A�OZ������a��.�|���nh�mh�8�n����(Ap�]�'-
q臊�X����G�S@���&{Ӽ�ΰr�o"�]LSGH��t�wK�$�2�*�c�`4��[�>Q��G��-&���!̠[~]�!�W��W�oi.�v�&-#�����#�Y�M���U�S�R!��r|�����_<��u��� j����M�0��J9��g����$���u�����t��2�g%�t�t�^�=B����������g�A��%K��?���YL��t���8fC� �N����p��Q��o��I����,g1>;/��Ob|r���8F�g0�|�%�F���ܓ�A;C�sj��͊�*04���5��z��e倪RF奤�2*��p�e�dx'�	Z��ۀk
n	�@������niG�� ��S�n��+硡e���\���X�DG9�\wQ�v7fW��|P:���rf<r9,[v�R�s�S�,�e�Ѹ�rNO�$`��1��p�t 
O!���!���48�G�-sUh�N��k��r ���M���K�4�����%�]3JWW�/��}&�6=8�̟�lSZ�Ne8�]�Oۡr�2�B�w#xm���h�^iR!�`���Ulz�9��t�!���S���]�^��O* +�b�"�fH��-��r�5+���z�5�ׁy}��=��^�=�&F�_+����S����u�/(+���kxRX�N�6��P%$,���;�* Y�(�G�tT�/���<�ٷ��/|�5M�"��%�I�7��c�kkz�*��`A>Ʉ��P� @�Q������c�C�9�\>��GU:�45�/1��!�5�T�Ju���t�	��wQ�妌�&�}:&��/��ͤ�;�)��2{���8[������cZ��&��K�4d���$e�i�9��|BE�4�ZoG�;szM/��"JJqs<���'L������i^mz�R^��\)ɟ�p|�R(ޙ�%BU,a�3:������ɶ�I�X��*�����O�8�[��Ǣ��� �򋨉�3��`���b��\�9c����yQ��A�a����X��0�������1{�q�����QL�qx����(��;Ob�g�c���AL�|�7���[���;w���;qL������������!eρ3�x0�V���$�etn X҆�:E�ԈϙRӒV�O����Ơ_C�T&�6D�LPt�G�e��c�I�-ey��%Yv��L����ކ�i2(F��na��^���x��P��`���1;<�^��l�bw#F�f�=_0��>�Ђ�U"9��;;W�0�Q�ޫ{׹�@Q
����{�?���7"ɾ8�ؒ���2�?#��"�8���X�kx�원8��C\,��s7Y�!5�D&��g�IMN<s�F��mt�_�] �}'BKVD`)(��=��L��rd;����(t��/V��C��N6�`�So09�k
0���q�MO<��.���ap�2@��n�� ����n~�Q6�%+�*���AgK������?��T4b�ø<e�]�cT�28��*��u6�����`��!���W�_�䠙�<��A��f�h�xP�h##\�{ٗ�'�R㓞F�pi��U���>ch��I�.ϣ�屘��)䑳�G�n=��,��Tq��{���BZNo�x�h6\����X-FI.��q��W!��-��eI7����ߒ�U���勣>�Q��/�Jh��Y�<ٳ\$b!�  ֔��Y X� �B����c�¿����_��Ro��}��R�����ê39/��ᱺ&si�*鸒q]]�ҁ���x5�n��NT����Ȁ�>�:�V�~~���NW��?�x�P�Z�	��o9��}�,oF�ӈ�gQy4���a�t�zØ=��yx�p��Q�Ɠ�E�lֺ(������U87��4C-ƣ�7��Z�d��|�1#(W���aL��G��?�ѓ�cm|����܇�����*�}��t���818&>`�w�ROH�x��_��Fg��+[q���Z��s��� gØ������G�G��Dt��V,��cҨc��vNqP����Ǯ��e�"Iw�ør��S?��g̰,��08��fdM�'?Q�Y��������t,�_,8��)Q(��i=�C9�����A��Ep�"m�)e���N�iA��Kt�_�ݳ�&��̬�Uu��bD]�1E9�P�f*��l�Ϧu/j�{�JN���rf����3Wr�>�C��?%��CQ`��>)c\V���XIVD�#�);=�緟ƣGOc��NT����|9*p�N�k���:��DT�ۺ
lh@'HIe�뱓K#��]N����1�'*g����#=<�+��ԫ=Rx�C�ئ���l7u9�M�ʬ���1}�ݘ=�F4.FאQ(�^B��8�Z{@H�|�>Om5[9�3��Ub�R�(=|3N��Z���fT�O��Ű6��T� � ,O0��eRQu���3d�Ō�4Iz�J_
R)|�����y)[���Wqē��c�J��t�x��tfTB��G�+�|@:���`�R����/�M�R��c�k��g�9����eۼwܧ,�,�4lH+��B��OX$�*����ٱ,�VI��0ri�Y#�B���+�����}���
����p\��(!|b,7,FN�g��Ս�䍝������+�
]I ������a��,p��Y��}k�_��`�F� �2��Γo��h�	C;%���J�^�����Oc���Q�F.E�	PЉ�?��2���O�c��oǓo��q����`���(�!��/k�P8F�aP����Bn�4zXe�ݢ�TxP�I;���t����V�v�b����1�|����o��Ө#yꍵho��um'(�~��,|�b�d@�E�s_��f|JzF�c۬Z�e�,�2�\2���m��� &q��*u�p������UL��@�4���v�8 ������sC�e/r�����X�� ��f�s �0��O����A��D�x����Fӝʢ�l�g@�K�E��5�7����݌N}��'�?���G1�?�����M�4� J���d{܅}���t�+�������u��^��~3�O�����TN�5w�Z�)����Ճ�þt���3���:iy��g� �7���N=no�r[���
Z��I`^/�J�U��҇��\+𲏩k��6�����Q��vt��0Q�����t�f��v���N]�3��˕����8��'Tu���~,ߍ��il̞F��0�|_���g���ey�d������)�e�Z��}�R�e�r(�I���c�/oj�ؒ4W�����r�dN1��.��=��҂�d�{�b^28�W�MNs�+��6�t��x�@��f�� �yYa��#��^UO"4q�O��?k�>�����e\������V�2��J�-ܠI�/��%Rfp�uD�I�*DȈXp�ڱ�N\6qɻ��9&^@�|�m,�[��s�����7�p;��/<��/�����X|�˛Q�� ݃�w�P([i�2h�����X\��W�>�y�sMb��r��F2�s�F��rnx�-�~=�|󿎣7�aL�� 9Dm���=���wA���o���v��������@x)�	v��LepC��d��(ZXk�F#6Z���m�N��d!�d3�](��U��؈ƕݸD����FC9r����Nbv��׆���v+�7�b�0�_��DDa@%2��}��E��#Ι7F�/�#�V��_
�dK�5���
�d4)�#�x��\���*399O��^���Y�8��6y��˭S1�_V���sd�l�A ���)Lh��<����������8�����4-o\�I�%���@��Pu	���[y=��x��^�܅�+�����N���"��]�A�V�����4�pE�CTO��Vܹ G�p�}��86+���<��͋xy}-v}1ۇZ��Wv:]�G����)4��K%RpB���GA����A襷(�^���rXJ�(O?��<Vu����w��>�RgO�W;�&
�9};6jwc�3���6FV�ߌ��\P�Z��) ��"�|��7�&�$끷����smWz�x���ӊ��oTc��g� �[B-Y�١���R��f�(-��/�Q9���]�7��#�y����~�~�����AI��l^��t��}��s%���w���3N:�6����?lLNs6/p[�6Y� ��#q�,�yQN��	ޮp/g�E1<W�}Y�\s�����&6y]����1~���u�>�����'1x<(�@�\�C�7�t<��>
¯%�UE͆�N�]��������>���݈�oV������������������h��}.^�j|����[���ǭ�y|���x�v=��Y��_n�럹{}+^|��[~�s?v��q��U��N�v�vO&W ]�ǜ��;j�͓A�+f(�����hm����@d-��?'|`~��2#�O�� 葷�}%��/�!8��M��ao1�G��(�m�7�ڱ��B�'�h? �;GC���k�۫�r�4�i�_��� țx8'�
)��nצ���je��ހ�2����"�n��ފ�+�1Ci���E�y���G ���#� \Mw	�0�B6Y<�*��խ���	B�l4��)��(4��tG��6�A��F�U-.K����x�G���e�|0��<���B��ὖ�N�wc�2�:� �6���kX���8<����;��]�m��ֶ{���Ћs���z�/��q�}�g�+x<�o�4N���h�F�pc��z7�1.)�"v�
���'��P��%��*�O8����>tz��EۍJl]�x�|֊ܨ��սf<�����T���~�d��P��_⯐�Uw�f�4t6�`8�^W����F�gU�JѤ�K!�*�Ux�_~����ͬ�:�+sGE9}��Jg�Mx=��)�2���^Eѭ`zO�⫱�8������5<d�H_����+�cV߈�i%�E�,`TYd���m�:�qB�YuIO�����z���#�d�e��y�KPK�yd]�L+a� O���L�k�ܞU����8���7N���ĉJ��<T.�qK��Y]ƭ��?���r_1�����Z\`�\�i�$�VS��'�
���x������A?���|��@����<<O��{�3��ڍ��я�����|��<~�����b�r}'^�x�����ӈ����p;�h����D�	������k/����o_�������/�H���������M�]D���y-:�q�l"�f1d��R�A;�F�����f��]��WbWa\?� �%���$R��N�m���ըn\�E���ۑP� �z��l�8rg �����U9���SA�� �A���C��!�2��q��-�%���j��20Pr����:Y]�����i�e˲���*��@1�nƴY���(l��F��L�T>�f��pU �9���lT��"��O~�hx6A�P>�,���Z��'�@�0軭�VT����k�Q3�?���4Zb�}��
sN*n��3ux�!+f�+���P�n��۱h_�yk/�N]1�>>��G���\�e�ɓ���/�����d�Z~j�2pK%�֋�F�!�f
; &��fi(P ��Y��c�)O�́�1��f/�p�|Ʊ~-����d��U��b{�j/���p��)
�F���L�C�*�׻p��-�T��&�6cQ��Zw7��f�/�p�E��\�^d"����X) I*z��m��e�\��ҝ.z(��l�1����[����u������@N�-�z�@<�ok�E�"mx�Ҁg1BZ[��q<��!F�%��/�*x���K\��F�*>FL�)��0��'��9���,���-��o����f�;N̔u	D��\�	nuX_Fd$�$�}'<��^�+���g
�S[,�����jB��$�E���r�����3G��/�I���!o��R�xC~��a�L��n��SM���?�΋38�_E�����;�S�XƕC�K��tp'΅�pPR�v7�>����/|!~��Wɇe��{[{q���/s��E�O��������û�ۜ��N=~��C�	�=_k�c��͸v�ŸAh4[ 9�������~�6��r;�{q�֊s�|��=��5�Pp�v-K����_���u�i3�\����H$���d���nԶ�c����`���dI�<��NIIL�a;[!TE�\���~?�%���VZ���j$�lv���=(_(s9���WX+[t���l��n�_ԕ�V�e��r���q}��6�4`Ϭ�c ӈS��)^^ ���)
�V��`����ù�:s��� ~�E?R� ��P�5�NJ6��@Ѫ;�i��,���}�� �;��j:�G��a� ]�ӈ��:��w�����*�|n4Q�biAG�,�ݍ9�I�w#�խ�4ҩ�Jz�H~WHڮ\!v���v	��}Ҏ>^� ��Q%u�ϕN/ ~<���Mk(�5=HD�����x>��"�bvz��<�8g�܊K���y'�r���W�4��yo��g�P�z
O)H|��`^��tv5�+�ry89/�-�������:ʭ`+���ǚ��T<�O���i�2u��y�ԛ�
�1�Pl�֍�V��]�EN23-M�w��\��
l*�ӓV���Jt|�k@�L���5��8A�1v��M& �8 ��ȶ,�!�xl���ad��i:i�	Cz.�e�ɟ�"���٬���RY ���'�d6�A���<;��l�We���ȕ}@�jz1�(w*�1P��\�ץM2`��_N���p�b0&�_�ذ,�
��He�e��2|o�o��:��gD,�l�<��a�V:(=�o�?�����ŋ��J�/b�W��~se�b��>s�?�/ƿ���.��H8�
+ğ~�;q���x��q��i����
l'�a���G� ����	�t����Jn��r���W��F/��;���o��^������Z7�~�FT9��9�B`9
i�lm����ӵ��Ĕpd��p��lRبVo���*(��
L&��*�}�0������p��s��@�U�L�[��-�F�L�CK�W����s����w��JY���%�v����h�x<���(�Xŕ��;�^)ss��k.�z��皞M���2�1ap����ׂ�d,�c]
�Ag|K��p�[�1����� 6#0]���!.�ܳ����p2��Q&��@_6���v;x�<M�63<+�!��j�1�gл��[��u<��1r�`ڨ�t���}<N�qs�W���^���%J��R�~�R��@ht�ж��u�O=|�>�D1tr�{�+���lm����\x%}�2^�����~<l��r�>�t��:E���������5U��0^�{�� �Q�N)ۙ�|g�:J��rv!y�-w�Ww.=k[R@���6q��G9��qS2�&���x�A_-:����������i��-q3 B0y�OB��#������lU�b3���dt؀2�.�"�@�	R�9}�L�4ߑ��64�H�7�Z����"����:
��!��2��|�D>�/}n�I��?��_�H��l{^��_5Hya���_94c䱕QYp$��\���eed�u�%Ⴃ㓈�V�3M���\��1�uz{˼z895�=�V�:���8�d�Ľ�c�lPX����`��.�Ņ��Tj>���J����;�(
߅�]�Jc3�\������&�N>���z�S�D�oh��{�����` �@�f�4����?�ӷ�?������}#��f��l���G�9n>�|��t'xS�w����1sJK���i������k/��@W� hiO�
	��4Y�A^���-��7�s���	�b�8W/��s�J��v;}�cyɘD�H�(-ӚV��q�@�Q�Bжv6bm{=f�ՇҶ�r8���(�x�B��T`	�f(�͵���2x��)m���a̬;�S��M�U�R�,a9(efa_ҷc�)���N��Q�&��`*�j��C��m��1�C?�Ԡ�om���Ju:SE�uze�Y�%��(��.�D�M�שOQ�����ゃ��-Ȝ"@8[��\$���	���>�Ms1TXK���CM�t��?1�pHr g��ǥ���{ۙ�vRQ!�A��|����#x�f����W���S�5�����ƨ Ȟ�Ǿ,���q�.]��}]��n�!c��Ԡ��0��"��m�+3:��yg�A�v1�V=�n���,�r�o��eҔ�q ���X�����|F?��$��`�R\�6���N���z�~�r��vk���p�Θ�A��ȿ�r��ъמߍO��76]杤���Ki�G���r]x��a���뢨�Zr�p�{��d�:S����~2�^�dQ<�:�ԙ��?��R�,�(������ Âr�i;=�M��q�ٚ�����q�_%�*����a������:��t�L��ȸ�T�f!�k���h�1`�<ͻ`x �x��y�n�r�0TTx��0.�'�_�ѓ~�q:���q<���|���q?������_}��߉�����������ʫDog+n��Bl\ى&��-G`W���G�
����J�@w�6���ը�����p�+8˲G��|�0���t�5�U�g��y���q%ٔ�ղg�i�&3�`��QX@Jf,�L!E;� �sa�WP@��G������	���Va< �z*�%�5�ϗJU�������HW�G��:]w��f~������h���s5��W�w�ـ�lw����sz�r+��H�� ��N���sz����~�P�4'x#���������*���<� �J����4�
Q���+�/����o�G{�w�C|(�B��rg���!�'��S#Ds���y�I��\�H��HS8�_N��9��,��I�pՊt�K��r<z,�۳i6��ʢn"���x_̥5�4Ĩ�v�v�B͞<m]n���o؄����q1E�=�E��&�����l�m��S���f@�|>S3�tj�ku�g�0�l�&�ouP8�ay�H��d���=��_�mGc��~?��Mi�b�B=�Y�>Ex� �+�h���A�4_.-��4Rǭ�,��kćo��ƺ��J�.UF�+���(4��c%x���1�i��O��U�Ȕr��^-���˛T4)��<v"��PI���/m�.c�y� ̞�!�U2w��˒���[�BB�̟�5�d������e .q�_��	�\{������*��L��� �V���ݎ֥�8OON�t�S�f�޾{?��Oމ?������޽w������ş~����A��ϱJ�1@�������B�����i}p�l���b�g��N�t��/&��s�Z�*&?�����T��uN?J������qp���^�Lʠ5N��c�9�l�4�r��_
:�w�v��Y�� #ZC��5���.�.��wq�+�k~��ۆ�U�#\�Lp^��_d�]e �N"���FH3���H�ٯ��L�#��I��W����Y�$K汄�j�
�O�ǤvJ��M���|��yQg֛�aQB��C�S����p���Da�;A��h_Q�ބ�8�PO&���"�#�<a@���LW�g tܻkk��?�^�:G#)*���w�j�)"�ˤ1NUO]��4�(y�}��W(�w_Q9A�k���$�;wV�$�7��ռz�:��,B�s3�
��$.��"<��\.��N?P���3JO��j�)ԩ_e�W�ƘSK����G��
gM�Q��9��RCA���6��K�(y��.	J(J�-�Ϋ%��	�����ڭ����S%:��+�e��e>pJ�$���8���~��r��_\D#���\�{��Q�]�zn��8��PH������n֒3zˆ�[![�`>���.�y��ˬ%d�P����X/�
�̓�F>;�6S����B�u�Q,C.ֶ��Q�(�g�:��R��r������/�6	��	��-����.e���9q���GJE��_c
r�͙��J�#�� ڏ?{t_}��Q��L��7���1�8���{�8��=�w���x��oǣ���8*�a�u�+���K��S?t5~�^���~%�OO���S "�@v4���iTFӨ'��O�h����[(N��9��=�JOeC�ˈ0&��-M\i2pr�6F߄�ʳ" @��e��Ғ�As�:� �����i�4:�'|'��禀�{�n�t"g�g݇�G�,s�f]!Sk�z�
���1�B=�V�S��B��t�i��~>{������,>T��E9#��N��]8��T���rez�&��s�2�t�3�P�h�gQO��)8��{]2
+�A�3�X�Z�Mh딑JI��@���ޙ���o��мڤ]�Ȥx`�hy����M�Qpu;ո�׉�W{�w�SF��,�U���s��=��N�@UBy��:2���e\�t�l�WIo�i �p�*&��?-x��<9y4j��L�~^
'x9�
�8���I��r��F[��[�;���wz����˺*���M�ؙQ�NǒN��.�	C�*��ě3a��\��?���z�>u�c�l�ĸ`̺_��|�,۔+��:�T��ƚ��y�Pf.�iu��ɊR[l������h�s�8N���h��uм><���Ӌ��~���u�z ��ۯ�˱�E�Xs��t
o��-��*�Q"R�#��3%�y��^�Y/����y=h���,�<>�� *t��e��ܑiD ��&Z��?OIO��/�\M�j��+������rX�{��������������xp&Tj�o&���8��P(niA�s��~#�G�G��I�}��'����w�_�Y<z�N��3����'�'_�gqt��tr��qr<�"iĕ�Nt�`��Չ��z�_���!����;��~p�4��?�ø��8<_��	L������BX�4@�����IF�����Q�J� �*ZPD��� ,�X���&�D�>�l�h�\դ��A��O+�k�ȓ���!�K�(;T�	[�<J#`��.*�ÅSM�\��� !�S�[1o��`��sy4�:¨Q7�/��TN6���S����|F�l:�f���q{4H�p9 �2(�6�`������X�z��<��'�i2Z�U�z; l���K�F\0�sSGP��Ձ����}\]�XaS��Y�	S��
1�ae�	�����!���"
_�9@�_�(��Z�$�Ge��V<����"��ra�KCŁ{�eN�4+�#�.��Cɰ�w���Rc�"����~-{Z���{uq�h�ϣ��P�>���\�	#����R�~v�6�p䳼i �x��4�����4_���l��RǙ�p!�^W�h��8Q���$9��4�3D̍k[�[oR/��|���T��L�g�����u����/lN����S��*��V.��x�9����H��������/}����?G
]�ٜ�!�-YBid��3P�>��x�͗Sh�c%�jK�PG��|^	1�ܦzmNE1�z����<��XE��b�۶l_������K�� e��3��J����a��K����>���ۊ�t�K���t�o?���I���'�m]�ǰ�`-�9{���q��wߌ�������g�1�SF]P�3�#��k�n��M�J#6���N5..Fqvz�Ǉ4�؆�o�֫��k�>?��O�~���7ߌ�{_�?��A\��Ѻ~-f0|+ܲFh6�y{���.�E����4�e��*7�6�k��"�����4<c$��Ȕ֪��de��5K2
��fo��p�{�Nw5�-�'s�JQ�Z����h��g�1��(��P�i?�]���n�e���^D��q�{͋	�%���&׾���%Jl%�L�;�qA��磘<>͏�5����CH�d
��>�@�;1��I�j�J/:�vs����4Ο���������f>4���Ji�s�����.�F���8Ǔ�����$.�z��S�%�v'��[W��,�x��عY��>��E�l/<g|yO�کĕiQ�wZD�����_�9X����P�Us�3n��s�i�$:g�K��{��r$#�W��@�He��u*=+��98�c9����,!$�(�v:3���x/Y_�Ϲw��� �<���o�7�
�07�x��O�%����p\�.�/"L��pk@�f򢴣}䐷�V�+wDh*m���9]fs��.���['�_�Z9��9-�5
D?�c �gz�2�O%��ĵ�t��=�\!��iU�
C���q�<fL\�j;���Ib��v6��;�,�2����'�g��3N�8����?�|�<�%{iM9J�m/�C�K��+�/�R�����5�ęH������q��>�w��J�%�ɫ\,�;e\1徔d����)�r@4
;��\���x>���_9�~����,�+�������J�G�������8��ߌ˃o�Ύ ���	E���vXmm7:;(���������z��x-�V
g�U�Z3f#
h2��Gq�[��_�V�y���ps�z��z<\�dc���d����!��#�?�)�w1��h���	��p�؈���3_�x�G��添
�qُ�X�7vt�!��bʶ�`�p� ަ�N�B+�*�!��k�e�����W��A~�!&�=u*����GU����Se�Է7�6.�;��?F�o��m*Y�����uF���ɾ�@�6��B��r?47k]C:%#ˠ� a.p�6�A�B�b���ʤGR�p<�1���U��V5b*���p(g�s��VA߄�k����|F��7l&�'Q�3m�	kN�m��L��R�)��/�x9X�/�����·�ԛ������/_��s�F<�����ȏ(�i~�4�Zi���RrU��9�@\
U��Cj��8�8{��8��Og�'���#�൸����(ۙyT"X��mȏf�����	Ц�oYa����۬ˈ,#\�iմ��A�9 ���L�����zZ�zW'N��q�w� t��j����OZ��W��ƙP�Y	W͎�9�<)L�A �'�Kx3����]��mp5l�;��fa��Qj��E�	QLP
���Ȼ�
ݜRM��J��	�#�����H�UAϑ�t�/yD˾Me�%K�?�$�L�!inE,�����.�L<<��۱�ɥ���*�|)���#yۋ4��?gL6�2�j���)��
˞�-���(�PV>J��?�rT�����_9<�7�{+޽�U�%�'���jv"��R���x�r�ɽX�����nk�V�/<+>��սݸ��y��۱��}u�W��i����m�E�U����twg�ׯm���NT���NNb<<�����T����X;�/ƮEa�}\*��%�c|~Ӄ��8܏��1B�%;�:0ϠU��4���|�(��x��>���蠸>���s�X��8�R���ҭ[pp�<5w���:V٭>|�4��	�g���/-�
�_�q}s��]���C�09��g\.uu
c���A�"�Jer��C�GMCY����l�m����pe�Q���S�X���vɻ���CO�������0y�Km�9��ف~�e��k�s����Uyx&�"@F=��g����"-�5<�^%��S��Q���Өxo�N�h{c+
xNÁl]]�F? �{��CĠ��nY��"DX�"����G^�V7�K�	Rz��0�O����r��������ˠ����RX��A��e1�'�H����-R�Ȣ��I�
���4"\ a{[*O*q��	+�G9�s�<�7 �aG����R��K_��\�@�����������sA�o~B<��ʆf�� �%��a\�b����J��R��k7�'o��vIW���E�E�`��8̗�Ƀ_Ng(���gW62Eo�nW��)���v<��XglYG
VꙌ\�*�}1��X(~���7��c|˳������j���il�JҤ���y$m�eV���D�<N����4�0T��.j�V�@��=T�4VN\�2���L�Y7�
�7�7WI�g�!NyCC����GA�RW⓭,����ʺ7�B}�s�!�SՎG��&���8AkG��-��L"��5�cڪ��s)`V�C�8?���+������6^M%���Q��t*����C����UB�n��,�z=:�|�`T��������q����!pt��P|���'q����8G �N�A���܃�2��C(��Q�.�cv~�}�~�`�Pf�gh��qT�)�h�����9�N��tHY����#,{H��ʺ*B��k����)�6�1F�AX��֠]��|�+�˷����.���(��Ad��s�H���)#НtY��n�q��Nq��ĥ�1��&�dF{���)X�Z��nE�~i�E��"\�\���Tx$Y�mtp��NM�,���;;-�grY;ޯ�~�g��f�*�7���DY�呟v��݊�,���B��ҳ��"��:�+��,�"τ?����\&�9� �7ާ'N�K�+�|^/��o�&] ������%0����|�"�,��.a�X1j!*x"/}��"HZ������R�<�v�j�#�=
x�(Or�2���Vp�gL[��mg�!⋯ ��x�}�X��jX���¢�ǔ�C����!<�9���N�_�gCw<S�S��[����huʻ�@B�#�¿�,�]���(��!p����ʢ�Y�/G@֡��:�cKz�!�A!M�f=��+^���윟���+ �-��BA"k�gV`>�?
6�;�󐇞�1�� �K�/0~�я�/>U���2�彁�<�C0�H�y�����[�9yF�O�ee?��0,��Š��Ѿ�BL���{�g�ҋ���5�t�%>��a*���AW�([�>��%`�5j\��1@#��ബ�C|����ZޙG�T��5J�|�TZi�~f�P����������G?Ͻ�jN�t�[(�=��g�����Bm�?��n������;�w��N�O3k��l�~Gd\6���Um�<���q��Q,�Q�1��o��!��0i����0�+��њƕ�e������6>���>ϓ����tG�v0��0���Y�}�Q.Ŕ�e�H<[�!��N�#\��tªS�0_,�Ȏ���� �,�K�S��-�Q�p�O���u���u`�2�8d�9���:M����O{�e(�39ݥ�IEµ��q\��|��%͙�:�;�[�3_�1O�%�,K�3��Q���)8�K��a���
*��n�݊Vpa��p
��g�sJm:�.c"^��.`@[I�E�/i�������	����KA�F�/�PrY�ޣ�ĥ � px�WT0�Z�8��  �ć>�[�EڄK>�^�_��kИ����@��ﰜ���*�)}��!��?S��1�r�Pτ��|L��砵�Ǿ�q�;�ȧ�S��J4�����2<��
�4p��/�"��4�˚幥�W�3�b'�,]}=C�z|��]M��z�m�*N���I�r�>7P��ƃ��8u����j�5��Ճ̈�=�( �8֤��\���D[�����vl��T=��m�2qK�6����ք��Q�T��������i�c���w����r|��d�=��0F՘�6�m�[�*�-�쉺����R�d��[*r�GN�i�c�S�xO��/�xk�'RF)����@�<��|�Z��|I7aZN+\G�U	I�DB���-�-Q�H'z�m��m>�@��3ጐײu��Ǐ���!�э��z�)�:����@c��"���0�n�=��r�Ռ6B�=ܚ=
f�Ո�Jm{37s���Λo�ӷ��s9Ĵq��D�`�0��\݊��v�7�(ы����G�'��i|��F|��q�\�!:�4�'�)���b8�)���E��1h���Wß�,I�Ys҆�����R��Ђ�5a4����t��Ӓ�v��t���Z�Sh��])�T�r���UL����3RƾΘ�����fr��r�p����s; ҵYW�3�L	.�,��d�t�Wi  �>6���z�c���g��.�����89<�]o�� -H�K>��Ϯ�W�)�B"������s'�r� �ڝ2 �\��T:���j~�ԗ�[~E��\�oSr�"hr��VrnW�0�]��_g�_ɮ#䳡����,��H���g�_l��W+Q>�g²��,N�y ���@}
�b�'TA �3��ŏYB��ۈҜ�Zc-6}���*Ө<����w�_�.��x
���CXe�'9��o_\B���ń�_���d8`JyS\�8Rِ�2(�	�;E��g˯��| �B�Uw�ʲ����6� ��w	���o'� ���sp�������rJ���u�>0�nv�d�7�����)Tx��g���"7M��I��{�� �c�QR~~�ςW���yp�����kʹaqZ�ZNU�� ׅvrG�6�{o��RM9����/q)�R��<����j�4����IR:+���O%�h����8�ڨò���ZǬ(�i	���������W�ϧ�w���y�A��T�E���)7��G�������0���qG�O�!���.��N�G�`��׶=Ci1iZ� :��ڠ���`�|g�M(]�p�/Q�����M���]����x�V/�[�ۮĭ�v\�����V�[��6�7_؍�|��x�c����0��0!����V/���|�T�_�� �zITZ�
�B��w`�K�s���p���ʒ�w��MA�`��ǹpb|vJp�e.���'�VԶ���'�&N�� @�cH�
-
����Gp}q�ݛ�F'�>�i��!�==a}��F��#	@����YYK����F� k�U�"��U��(�� �N��`W��`լ��k���ы1��e9�vyx�S�U�J���� PP�(S1���;O��L�ԃ�ҧ�DF:��B���K�*g�To*�2%���L(�b��%L���$G�B�����I+蛄�Hb�%&�tp��X�����g!�(�Y�qJD*�~O^�sy��'3���D,�<_��ZZ8Mݣ[��o���#a��Hc�(3�p�. �]}��s�p+A�;�K��{`���<�
��@W$���1����C/'m54R���*����Q����]�����5p괭�J:b�Oނ��{��F���;yrJ����g(��#dM�tS��)����0(�<bGڿ�qJ��[��Ύ^�ۗD�����!�O�甇l�by�	~��b�]��J�g�_V�B/������/e���ƅQ�O�U�
��#3���JL^��� �8-o��9��S�K��s�K��Iy"��%0!���)���i�e�Q�?~�$~���F����hf��<�o�ㅫ�xx�(v����>R��x��7�����Z��������ZĹZE%B��iAӎ�Ҵ�!�NFX�C<�+�С�\I5�Q"M*0U�Ʒ��U>�]�Fl�!}��f|��-�ҏ����۱��!��I�7�]�O�����ى���}��?������x<��˯<��^�~}=��n�I${�>�g<@ږ\NGq�^݂�U��P�z��Ѫ6seҘ���8QFg�iM��o�v�A���)J�<�����
�`��vt_��n;���<!��'Q= 
D'��o��x�	Z����ڊʕ�8�óQ\�?��ݓX�%9�R-��
���Tf����X��+7w�����6���������h;&�ɠ�pQW]�����u�慛�_o�9x��1{�a��#*!s-:�T�=wo�TP2.�e|n.����s0p��$��8�}�弽��"�C�"/�M�ʒ2�yC� W"�W�0?_`%˷(]�9E|�L@>Ϸȩ��U�)�zLw��Ux�¶@Z�G��C�e*���6&���xsչ������Y�z����^m�mW�>�m6�9�>B��E��C-n��,.9WO$T@��KТ�J�b��C�OO=������8��/)�'�UdRY�f�%~�WN��\M^Κ��q�r*�4��-/����?Yob�5�	}c���i!+�7���XR���T0�G�}�7�!�o_�ى��nTZ]�(�	�>&���������NO�~��^�қ����ԭ픟�&~�6wE+��uq�F�޻/��0�����tYK�i_IH�%�7��"���Vƛ`��koӐ�0��[V5��O�����H�,�q0H7���L�x��l���r�@i$�d0ʥ�l#q++����'x=����Ob���B4 v���q�J+������d�4j��x�����	)�N�%�5PB�d�ܶ��t��T��ɜZsZCʊ��zǝ���`���x��1�5�ޟ�
m�Ie���2w7����l5�#����󻹙���9���ĭ݉ݫ{���^����/�s����[�������o=�?xc7�.6?�b����A0�����-X$\ F��1:8��/XA`�-c�jsΕ��k{0r�x�ا����({�ynKM�8�h(	���z:�ظ��݊�V#��1~|�wD��B�/����� j�Ǆ|@/�3HZ����9�s�<;��>8�?a02 h���|1�i�v��t@��2 �W�^�޷�ۛ�m�=���ԏ��O9���?ߗp.����E��@ חn�jH?OhG|�A��90e�T��TZ�&AxBa�S�v�#�.�n���g��(�6N'���3�x��#�h���L�֐w,Ŵ@s%���-�뵍��4:D�M�H�e���?)�J���`���'�Ɗ\��)��yLA=�
�;{�4>���6�9��Y�"�SrS�����sJ�����v���(@�Q��|�-9��=�ĕE.�� _*8i�Y�4��P&�F�����W¢�>��ö�q����0Q�S��yE�[)�u�3�m͙�LL(��cj���\��a	�z��x�zT�]�'���Ib��},0�����ә�ܫW7���s��Icdh���;6��Q�|���)Y�j��W!���<�C���	�[yi�`[Dm��n S�J�[�06��;����˺�ΜB���I>.=��N���qK�O~��5 �0�k?���+����-7噴��X��+a-�)��1�遏DT>T*���lU"���/�徑�r�	�'w8�����Q�R�B�],��8��9>��,����1��*}���US��N̓�Y��dL#�0�u�9#�� rJ H�`�K�$�W���-w4F��t��r�V�H'�F�!������O���^Y?.���>�o�)��խݍx��xk�go���{O�ǃ�y��]��/bB(��t��T�';A$���x�O����1p��Q,"�������)�9��nT}WG��l�7�c�-ǣ�X{ڏ�1
iX�������KZ�9٢bZ���V���r�O������K��0���kݘ�|��y���F�ۭ0�&
�S�=֓e�ʸ��.��v�8�!7�}�0o�b���z'_�]b~؏�1L�@��+��_��S�̀t�v���'����X��� �� 
����Z��@����p�����=��}%��X1���)�!uZf@Y��0��|�{M��M���=3:~�E�'�ON�ϭ��^H�&F@kz�;j�ˁ�ad���gy~VX�
+�oyN���>3s*ƍ�4��F�����������QU�u��w���9
��EΧb�@��S��������'��x@�
m�he�SZR���g�����9�_\1J}���{�c��A���;WI	�]}���q�<u��H��?��w�Lz��~-9��>�_��p5�N(C{֎8��-�>�[k���|���Sa�-6���z��'���<����|���(<�z�ݫ[������^;�m�<Q!泰X<��x�?d'�S� �ޥK�}�S�h����Ͻ�����?�u�\�0�F�
� ��ul��Y*^y2˚��*S��_�Y�/,��� ����D|��\�HT1��WB.97�42*��\�19e����2$ѳB���Գ����(�w�/��}�^~L.�<r~��h�֋�q�����R������a�>�Բt��F<?�HE2���XP�A� � 0UL�2>�H��C�� v��dŠ��c�C���lрF�iԹ��!��s�ѣ�i���� ������ً]�ս����6�#x�w���[XB��8�X���M}�r�\�Vŀ���n���T�j�$�o���B�OY������p���~{�A���` ��0C����2��k�e�+}!���%��F-j=�:E_;����Q�GT8���nl�_؄[}�6D�&�`�Y��9�*���}� Q�8��Я@{�+��\Z*��(x�
�4�֡w#f�v�W\�xP��(2>H�c��9]�f)|s� $�>�=�hn�b��Y�O�D��IO�
b0�}��peP2	8��6��xj|���%��,�O����cA���Z��j�.ȇ��>xO�s�6��2�_5S)��Qq�X�����i�:)6�1�2v#�2�"��i�������H�jy���_֓������Ę(Ɔ\�;&�S�t�<���r�<۟ߚB���+�x��s�	ζI�/_��*��I�S�CK�@תb��t8gy���2Y;�|?s]!T�����<p���4���}��1�}��Ⱥ����;dGT����<��W3���s��r٢�1���z�i��QԎ�6���)�1��/�u��\(�\�^�,�M)�f�@yU�[ѹً�N�a����4fo?$�]�N�e{�+���v=�W�s��M;]�q��V��^C�E��y*H ���脜�d��H�iA�:�n�|�榯�\�z��mSC�����},�gNȮ�p�:�r�Qwv�2�K�0�P&y���S	:��/���))Bi�'(���"��ߠ�C��UuT�0����s�B��D7o�{�%�8��\́q^��_�կ��E��o>��ۮ8�q��P�ʍ'����\�����O���I4;��m������\��&D�nGw�Jl_����o2X{�����c{w/z��۴Y��Yvp�Ѯ�!�G0b��I2��G�	�[�A��]��X��O8��yL�gZ4��V;^A��;}%�;.�Ntt%����^���mؠ�M�
b�~�:	���~:
�O霉��)�ս���E��C��2�9%���L#>��U<H[m�8ߍ�'��'x=s=������[:�N)MDg�P������U�جN�z�Ó��>:@)0��/;���u��/v���ѣ�F=v@����%�:�68���k�P稅!hk��R	� ��q����0(Q1����(j��t	;B����]e�B?�9M�����J�2>�r;^�ڈv�z]��὘#t�J~{q� A��W\ǔ�]DEք�syԇ��s�
=�Cut�K�\E|s��8���m��{���������K�=� :��hA�Vg��y�k��r�Z�د0^bL�f�W|�8�)b
����٣�T>R#V]�������>eg9aN����%�����	�.�$?�;#w@����Ү����>J!�M���ւV(�\���5�V8�G1�K�D�9A�"�+���)��[;���Y^nu+�j�OU�Cg��V5
,�4@5*�.���vܟ���<'�I����F+�z��3}(��W9e抷c�}�oѿo���?�qR��D�.�B����>�� m��&�q?g�Ր[��~����O��/��n0&7/���>�>�W�>J���)p�����VP��(�C�>}�Z\b7xU<�ݳ�{����Wvx6�N��l�2:����+C[�Mx�F�6�����^z=����\�A���1�z&iZʧ�) �,��g�D֬�0g��{w���;D���������:$㳽�n�Y2�p��I@�9�Z�{ xCy�O(����|�����}at�z{-6k4!ߞ�b�g|�$���1B�����������G�g�O}6^�ȇ�_����}�3��'?�~���'>�����+��/��_zI����A��"���'���Z�t�J��|�;2^+�����*0wfv)dӥ�X9�-�
�A�lעGO��R��L��zg=>�µx��ױ��w�n���v�uG	v,B""/������#���^��ǯ��ϼ���D����W?u;~����p�4~d{}��i�W��:vV=��6BƏL��������Z��n�s�Q\�b�5�k�~���V��g_�+W�q�I��P�:�Fk�n+F*��N/�ݺ�k�q��0��»6>�k�������+ѹJ��(�0��'e�R���t
`A���rx{�i����\���'�q����bc���p^���Bfm�����M����ڙ���<>��&}�7=���a� ����}�����vc�:���n��l`p���W7��_z5>�#4{s�Ǳ.�h� Q��~q3>�ɫ�/�}�F��8����J|6r�7_����Эj�*�q3-�6�ְ���we�����z=^��A�c�Çs�~[��]��M�(X�ɟz�����]"��\�i�K<x'7^u0ˋ�P�V�^�� S��\L��|��}�PU�nǕ}.^}/~���G}�ck�@in�㕗6�#����k�خƉ���
��qԢ���yy/����k�vi�c����;�ѽ�!m'����G��Z�����ҟ����f<>:�����9�fĕ����[��݊����\{ G�q�[������~���+�ֿ_�����Y?���G�l�k�z��Ͼ�~��Xk h��|r�00���q4?�Z���>~�/�x����x�ޝO��Do_��b�{�?~3:��k�_zu/no��Ț��0�{W����������ظ����rn��_���7c�j�>�gN#�F�ޫ}�X+@�(��\W��;�t\��c���.}�>�7b8k�9�tފ�YM��x��@.�'|�����b���=xU�Gq0_�K�h@^)��>gg$X�D)������,[fY�2Ɩ-㕏����{��yrr
���ix�?+�O2�|~�+���;Ǔ���<��X+*�N��P�cֱnwX��Ә`M�����{1~��6>����?�blnoE��:�q�����E	P�F�W���;X?�(��?y�<�����i�{��7\�Ք�ր�ORk�V�:�8E0v��˟��|�G���#���T|�S��kz!��y�k/�[�Xxx=|�atz��v}7�xBo�{��gw�ܩ�su}_,��B~=3�6��`?�]uy�S:	+����җ^���_�����ʏ�_������xn���~4��q�t�f������?��������1D}�,�q/�Kys=��ص��/}<^��K^�fg-�����f%�^��-<�����܏��+�xr�0���۠��ߌ�7��'������7�<7&G����C��v�W���t3>����W~�K�?�Y�� ��>.�kq9E��x~�˯���_��xAv��^��ލ��86��nLr��x{���O�W�ֿ���+������t�3��������l��_�l��By���X��Q�D�1�ƤV�~�v���'��ş�혾��[ts#��J4v��ׯƿ��?�������?�Y�p���k4��W�˟�P��/�,�����'����cv��ъ��[��/���O~:>��x2�8�{�8H`1�溛�+׷��}����LZ�<�G�  �Le�c�FD��2�!�s/�FJ�%�qD�c$�K�/�usZP�	E�*W�P\��t���8M����*E�od}#���������_����+�-<��x�Z3��ÿ~�/�������?���_��#>��WSi|��Q���8�tc+~�/��ѿ����~������gq�}�㟃��O�x=~�����~8��O|>^�u%޻�4�y�)hc��̚�����?�����g�5�N�s/\���~,^��k���7�'?���7��?��#?����u����8����1�������������?���F���/��w��*c���#����_��~.��O�h�����]�Ug���狽������/<>�q�QPE�w�ӗ{Ͽp#^`��c/�/������w���{�����]"1�����H� ���3+.��> �|B?�B��������
v�Z%D�r��zc��׾��⩠x�U�FF��%�;1��m��uW���Mc2rv��8:ˠ��!�+���/NH)��`'��%r��0�rA�� *�/�}��]	*��FI�>�cS��.��oh&�!++���q�TÝ#(�.����I`+u�%���Ln����`��U��nl�n��:�Dyz��x�[_�7���������i<x��x����o5�����ѽ����8xp'��c�tDu�z�-v�UE�*$�^��6��(��ʼ�rp�v�����7��/���������k1�Ϳ���7��_���+���a�?�$ͮ*Qx����Ueeyo�����QK-o2�0��7f00�~f��=� BHBy�Rw�m�.�mVz���}���|��%������k�ͼ��k�=��s�����x���;�|�z��S=�X^Z��W����|��G��z��[h�]�V�RFh)�&JLK���t��Y�K���Y���4�c;������hj-���������߼�?�;�{p�֍عu3\eJ(V`�����p`�zl�4���~�%Y9	�5
��b��ex�e�)hR	tْD^�}�*6���B��{N��O��lؼ�`�|Ifb�J���:$�b�����i�V)����v���4����F��u�"Iל�*�:�Ӻl�P ��8"�5���z	�\�|����T��B@}h?��m��5�>�`8�l���r޶F!=p`'�k�h�şZ�`y.�z���G0�ПB�TO�� ��ϊP�W�Պ�~,Q,Uj�t���R�SS���!��(�?��;G�.ܽw7�޾�GG�3؇0�ё�����eᮬ樘Tl+�|�ʸ�(PA+�\��?4��C�!�/O�Y��&�dIc�)Y�Z�L0I.�A�Դi����+kV�2��2Շ���P�>�����M�g�<������R�̴1P���{[��0ȼļ>j�A��HҲ�ɫ�_ɮ~?�ݣIl�0޺;����u#T:i�GcT����OET��5����/f���C����h)nš��Fow7
-e�z4�&�eZ��W�*˥^�l7�)Z����u�H���ٻx�["o������o�覍T�z�K~W��2�S�t�5�@�|ua��A�����䣏���C�~h��7�����"8����,2�A5Z��8�	�L�T-�c���K}l�ר�x�ޚK%�tI�?k���Ι5�L�E���5'E\���#����S��ܢ�9�B&ArYE�8&����J�j���P�̨3�2ɐ�X']y�Q� c|ƴ˓T��7�M�2,����2�<[��&'`��`�\��k�|� X�}�b0�㷶h(��(���G�ѢPD��t�i�	h��i_z�^c�5�Xa���]2���%!�>�thb��8�����w������߿�?���������O��s|�#����/~����>�xbf�AW��5AU3�}67Ci3���JBY��cMAj�$�EM�`7p��!2�<��}�箻p��ؿe3�nو]F�}o�&
��{�n���,���Q|��O�[_{�GN�u�&�4C�������Ҝ��WWH}K���a�L������Z�]�é�[�ש-���@��ux)�5�Q�����@��(SZ&���P|ؽqvnڂD����B��2������NNavvWn����I,��(�X�i��=a�!�Űg� �َ�۶���h�B�M�זE�:@��*�7gVp���B lfHk*���AVE ��-�x�kś}�6nEG� b�ti����?�o�:���\��B���SaE#���C�"p��Qj��ع{;F�1M[�c��]�@�y�h?�o^� ����'p��\��Db�%�}�1�t�@a�4�O�z��i�&lB_*i��"���ߘ^����q�VO����&D��\䳈ۇ��N�ߺ��\��F��o��z;���ie{}l'/\���E�4)��] ^$�n%֠	5���t��<K��@~1-�j�ua5�/l�#��*��ʷy�/��F�iȪGM��W��I����)*~��^
#�w����bUs��F|6�%G~YőK7Y&�2$*�0�����|Wl7�xp����H��2�u���dyN.��蕛�53O�YB��|�M�Ң�;�l�Fֱ4�2=?���f�'�^­�)��r	�<z+ssT�($���v!�~:i�j�b�wm��,���G����#�S�o>|��|���@���"�d�tG0BKxCW;	B��w<x ۶lA$Ԥ�@�6ʌL1���R�*:b�\���|i��h/��rs��J�
o�)���[B�7���M��V�0��f�&�]�Ϝ]Pu��|N��n���&A���쓠�+�7�Dʷ�4w�u����h4!��y��'�Q�k������\J�V �dH��PS'�BC�´�7�i�c,�WT:kuÞ��H�ӥ��y�X�Ν۟�+�u}�x9�I�3�HS�S�J��fAO��x����1I�P��j���<�,4ѫ�����sx���q��1ܼ~.�Ĺ�p��y;v/��2N�|�O��ĵ���3T���
Z�n�Vj;ޫP ֙�Ӣ�B�s�+�ؘu��eҟ53@��Ӛ���xj����§��6V4���fe��M-S�Y
�WN����G�z�s�iZ=�[(�Y��FmR[7h�ƹ�MӨ6�i��I��b��"4Pp\C��z���gP̖�����\�iܺt�'(�
e�v�>}�B&�'긔g(Z��`�����O������Ю���nLSۙ��cn*��Bu��A�&��5��:	�޶{vnǐ�2%R��~dɸ9*�+\��ŭ�Y�	�e�����H��������G�jȑh
�P�v-�H���q��-�� ����P��^:a��ڂ^�;�ox�A�>@�㞻q�޽�E������ή`i5���\y�A�7EҽL-�O�gh�Fl݊����䆡�P0���BWgi���b���'����FYR'�ӊ������{i�Xߋ��(A�C) K�_��3_�a�¨�T����d���Jj�
Z5�*�*V�o�Z,3���ޤ�ʯf�E��i�<2
����R�aϦY��G��Os�l�4�-1#��Da/	:͇�b��-8�w֍Ъ�E���r�F7'�q����pm
@��j�_�VcgK+뙯#B�o�D?�e��)�
�XY���N�#'09;�B4Zjx�s�4�B���<�8�#�ᥲ�̃n҃�e�<rubG�n _����o>�3�%Y,M�&|?v���Z��˧0>=�����%\�y�k�T�HCVFIc���D��"�$��T�d�uh	��o��t��:ZsX�G�1Ka�eXE*�T	@AȺaK�JsW$�����E
O�y��4��?z�� �G�$h���ndQ:K��J�Bق��e`��?�o����f��겍�,S��bijE�hQ�W*G"ՁDW':�0%)S���}�������pZ�")�0+26�<&޽�˚1�Qţ�m�؜��L�����@��a]�ɹ��z�����YA��O�V��P�7��L=�ݱq�bP&���Sp�Q� ��<�P�^'s�:~gϟ5�l1\iC:2�u)S�5PF!S@��%G �f)�)�lEj�Z���"'jB�m����
c��he�b�QzI�f��5�Rv��,��,/�a��\�.`ei
K���f��4�gQ���ҕS(ߺD&S��JQd�Z�`�a�hح�X� ��m?�H^kn�D��#�\���<��"��2d�\z�,�n����ޠp�>��\���p��E��p� �-�4�5�)���[Z��z�"BI�bm���p�05͘�
t�¬��?0��V��ZD�BVe�M�R	���Q��B+�"5���iLN�����
��@К)�U$�Q�7(|�|�Պ�F�{G����V5lZ�Ĳ���1�R�-2vk��ʛf~V��e�D /ih:�R%��+Y�)ܫ��eY�(L�.�M.���Zx�4+�*YR�	�d2�752ˋ(5��y}�;���=��-t���K��)��0�-���H�2�H�U��X�i}��Զ���#<j"��3\]�a%������c��@e�|h�@��E�pgC�q�űa]�f/6?0��oZ�{�6�]���h�,N�6{�@������{0�3�����ڃ��<���q� 6m���H76l�e�%�d����ܙ�B���I<u�J���aܻ� F�6S/�D��
�IS��_��"ˡN�p%SS���	�j�6a�z��D�����YZ&ٕJ����T���^Cuz�t`x�5��Q�WPѰp��uR�S�M*��X�h�u����rwc|�ՍuL�T�MC��˘[�>	�T�x_+fwS��x�,:/�h)�$����1<��	�r��)�_e��O�%�Y���7-�Zo��_:�����W>��c��o�.�G��@�,"�4�c�7�M�����2ٸ}�wctC7:���S9�o���+�rG�2��K~��bޕ�uH����i��-�b�7�(�2G�)|O����
_��r"�i����u�����Ľ��?��w��~�.���ލ��W�������s~���g~�����O=��nrF�ea�O�f�K�Q^�y9�k�m8�=���G �6i��L>˫�)w8��#��q�y~�W?��+�Y|���i��Ez'��`�z	�~ij��~�_ �����AK@�Z���<�i��y�y�$�j��'(����D<�MU��04�Z�RZd�hU��)���Bx��B)��H,���7Vے���O4ЛB�jqi��t�L�水����*��eL�L��٫8��	4��,(b�+�c-j�.
��'�5�T7���!�X��0c��!(����2j�f\��Ƭ7���������5>w�Ν��cW�qylզ�,�hɱ����&p��9�3+d̠ʋZ����q��uf���K���9ϼHCkb��(�ʠ"�SP_�Y���U��I�	�H��T;)��:�헰H:L������q
���������HD�!�ߜ�E�ңa�Le�#�#Qܳ��R4����疑Y.`��R����_��;I�K3����/S@�VɈԨ*!��x`s7�l��R6����7q��E\[�����.��(R>���Q�F}���/\ /��\�s"��� ��Cg2�b9K˒�3"Y]����jY��L2�y��Sf�&iK�Kk�E��?��A-�T����]��
��L�h-�Y!{:&�y��n�±ȲnV݈��gG?�ܹn��]�]80���{�ƻ��{�=����q��n��˸��Ә�|�^<|�o������a���>�ӏ�t��G�ľa�w��Xg��rf�`���]ط!E��2�\k.��0Ieb��:��6��۫2���-������A��!�®L��!�&UװLEirr�.����7�Nj́P3+E\�|�SWX5E ̒��c��mĮ!�4���S��p�QȖ��:#Hb	���q��Z�HW�d�rY~D6���F1��2Aޮ�ɫc�8q�.����("�1�%y����Ϗ!�
:��H����˔u�x|s��EY�e�9��_��g~Sg>���4r�Ρ�:�zu� �K�*G�r������'�Ƀ�8��m��=�$�V1��d���j.7�E N��ڣK�����<=�V{M���dU)�ڤO�$ZD�����3��!h����8���-��Ƕ�{;�_	ܷ5��[8�9�7�p�&��MA�3���֙0��څ͔�g��/R��R8�Lsɜ�A%�n�K�h�y�1���|N��>H�AYfM�lY�|ǆn38�������fIwB�\�]ŗ�O����G�� �v#A�0_.!R�!妰�e�-r�Z�,�<��gq��i�;�
��G�g��8���x��'q��Ǳ�{�{��� M�u�nKC��,*u�Ik�2;�,����3�´:tS{�0'��+
4)P�C�J(�0;5��񛘟����1�L\���(|�.a��E��pϽ�
&nޤF!!��}���|ܑ�}��x뾍��w�M�qWI_���53ٷ�rs��g���e��#�tM,��W���.���%dn�0Cs{��b"�����U�! ����}et�sck�D�ݚ�EV�[c����ʤ���j�^�� �1�|6W&�&-�ҡp�}�t3�0�OL�ʕ	\�>����^i`��F'�u����b�Z����v��H��1�BO̅r5���I�_�q�i�A�die���Go��!@%W�Z���4وi!��"5lIy�L4q��|�[/��%��|/]^�
�A3�#Hp]�s��8��&\�l�C�4���]o䑞����4����Wp�v2K��L���H���WI������U0i��$��a�/����Ӵ�/cbj�&O�|���8��l�"��h�f�Q-�0<�=;qh� �Y�q'��	c�(+y�V���&r	S�q�Ϡ�����^<Aa�{c
[�:���Ao�C��~K_���/���/�j�����c�?<X�������E\�v�o����)���আ��x��3���z�oӓ,
1��R�F�vQ�rcue��Ak��5<}�&����Fiy�٦�t�c�����-Z�s�¾�G�+��[��ٗD�����ùWq����YP��	�(o�GTg���(�}�,[u����®��j��v�4���������%�T=Ȫ?��y7'�4x'�'���}=���>XEoXk��#�p��<�_�<f����c����2�wS�H��x���R}]H��f���ي��BGY#]^�e���Jev�|��O�E�3Y)%K4�@v,���3Ykk���#�F<�a�6�����f=5�)I#;�l|���}`Gʏ8��k�eh	�?�e���Y���&��
c4�@O'��sHkޘv2���q��	Q���n�TGg��t���啠S���n|��1�^����:��>A|��f>�(i�����!4�3�p����׺l.[�syv�
bnrS�+���a߁{���|/z��س�s/�nۉ���޷�6o��ӁxG���iuNW�<N��d������,Z<,܆� �d�_J��P��m�I�/�C�hA,�M��D�Btu�2��_@f��K��-\�0��*��LHvc8�z@4G�y�DciE���A���]x��ؾ�������(��"ؚF8:�do�C��[O��-�ý�za��u�=����4��;Z�# hT��f��^E_G�T��"<�Ut���)X��՛�q��M\_�%j���=�Y�&H�WƐ��a����H��*2��~�/���+�8=9�ʟg��4@*��(��U��2��	!���hQ���s���0;~ϟ��6���KYL���
�Φ1��ʰ4��L�z�	`�h��hR��~n��gp��	<{�8nM,ba�Z�DnZ�)�%�Ӻ�'������.�Z��H�.2,iR_����u�O\� $ /qz��3�LM�5� 8�
�R�)����f&h��6!�a��O}7��c�f�������yb� p�#DV�J���ǲ���k��J#�QCW�F�a��'��α>ܢ"p��0��5v�μ�S'����s�QO������C!����˘����ɫ��QY"�.(���&����3�����%;�n����ɇs��i�<q'/MPX�/�f�p=z�D,�A�H���~� �����<��k��0-���-�Wp��y�pr�..��'��$�^�<L;�Bz.�@=?K-��:�Pf�I���u�4=v��{�<��Yܜ-b�R���U^ַ:�%��+n ��`�Sd��+R�<_��+�������2�&�	���-������I���
�j���0�UEw�Ja`��,��	�����+_���㬃勔���g�x'j�T����uG����$(w6��,�����dg��V������,b�����Pa!��f�N���i��z�<'-%�e�D�07 ���[��|C S�y�St0�7=�?��:lOҪ�_� ��ko�r�L��r�r��t��
��F���mX�|��Ǚr���|F%S�4���D/g�$q��6�(3><Wz)��4Pt������[9�����{)|>���s���n����k/ Op�U4GD�Y�4&�Y�#�����^�7��x������G֡�;	����S8��C�Z�<5���nݸ��WѬU��R�Zñ|h�(�WcK���m�]�@���M;o�'�Fj��)2�ᐖA��a5S�yTSL�`����,6����N�t�;��%l�H��^O���}���3]e\�8�K3GQh͠^E�����'�d����>o�Z�+�8�e�}�a�ۏ�2�  ��IDATM	FS.l�ta[�#3� �XH���>D����E�O6�J���R��36�Ǎ�2r,�l� �bKG=�µ	x�3(G|XM"�}�Ct��`e�Q�z}5,�Z]�ϳ��}�'����@��u���5Ɗ��k8��@�^75�<F�+H��fj_�)t2�͖m�85�E��)�g��e�א�@�7�2���:�h�������C� L���f-��r�B���֔}�f�:͓hv�0;B�#���B��Ao�ʐ���W-L @��*�W}��K�b=i�I����,^F<��VO���CAZ�ul�b �� �P�H+'�
�!�tQK�H��֑��!јD��A��W�U	���?��/<����*���n�8F�9���3'���#_�� �r�S-��j�Wm��B������]=���ÍK/���S�Gp��Wp����7�+/b��9���0�ٍȖ�0�
��
|Z����*���n ���:X?�,�T+����^F1�Bf�?�2w-^Gc�*-�[���0GŮ�C�'����뽧Q�2�G���>��}M��J��.�ɵ���r���<�D�=�iZ�s`\�A�5���r�C�?���4b���V�A�˃H9��2ǅ�L�u�qZ&� y��Q��� �fX[��,�� �'Qb�긑o�r��t��A�"eW}���z���u��$�)W<X�%�D)�#_�D���R�!�ŚH7�H��R�:;v��5�>֗�N
�:y>��^C��R��+ɬ6�8BZrW�~M��S	i�۟�G$���}KG��(J�p߁!��p�@ A
�"��ח�����̉y�����ṛ:_�ӧ'�����<F��6]#�8��*Q|���K�&5�I�m�[��Q^���֗�N�pB����E|���W��S�<��>,"��~�W?|e&�/_�FYs�:�"� �4�+UVt����gi=\��)زk����[��N��n�]O��?Cm��<�2�+�dM�ք���/�����
5���ϣ��l�ؒ�ZՕ��vAժ
Z�J��u�lh�UX�`!�iȵ
t�+���]芆��Ї"Q�%J���"��}��A�0������A�q��6�9��d���U���ׯ╉c�PSd����U�U�Qyoo����؏m�4F�q]�g��(v�&���Q|�;�Ó�b߮�U��p��B���0>���݃�{�6�ߍ-�)�jUj�XGp=��{���� >�wm��0ӹa*�B����T o�Սw?�ڊ����o���A�><�9�x�(���8���7v"H�o��x(�fgP��ȃ;�G����p��-�9�U�B'M�Qj�����^�ozx�v���B�Ap9B�R)H����=�7<to|�^��1��?-�6śx�(��G�c�-�NZ�Z�g}rݴ�Bx����>V�͸{�Fl�\��^l[׃�!����8�îl �c��1��oW��6o�҃'��j�`9o��O������}Q<����J��(���H�**�1�K��iG�.T�(���:��D�qD),��5twj5�a���cx�Vt�oBG�F�k^���!�уp$oKk{i�(
��e��K�"zR���������&�|p���7b��T�����u6�&P��{����ƞ�lX�j��+��n$��� o8���ڄ{�n�C�p�=1t��X���Qn�c�F�<�򦻌�d��$���<��ā�sw?^����0�� \�\Es�2�wă7�?���裒�R��Zӽ��$;�=��;���-x�ѻ���JRq�}Hi���H�k�Ѓ'����;@��F|/d�EF��R!�5qp�NlHa��^��~$�k[�4��EP��"_�F�G�	��nU�&X ���[Xh0Q[�-3_�}@#!W16U��-ZZ6ʜ:۝��*��v���]�gR�?v\{OV�d��\<��^�w��B"�(��^[�o��|�S���ӴZq�VC����"���k8��;=���y�5����|-�4[l⓯\�k��)�G�j	$(�:�ô	P�B�VztO'����jh���X�v8�?
�C*����#��ʇ>��k�|�|a�I#���.D�Ě`V��#�E[4��K(g��˹��Ǿ��¶��Л耗֋��t�:�=�g."��c�ΝHv�`zf.\����.���f���	�PT�I���,% i����d�e�C��&Ih�c�g�P'�a�A�фU������f�G�Z{ɀu�K�[�h�0�99,d��bc��@w2�C���E5�+P���+�c���2=Gk��t-ѲJѬ;��=�����t�'���Bc}#�<�1�7ڄȶaVJ-�⌮�[��B��(��zV���7�,P���M��C�Գ��7w3�����fp��k�ą����zc��X;��AP�'�d�����e��*��	>����3M�V�#�]�M*�折n�i�{p���ah7�OVg��C.���&�zkpU�q��m郛ë��6�n�㹕*�0i���b><B���t�G��]c���� �u]^<����؀�q

OVM�8[��2�I��|���0�ۺIZ�Z�����>���_�ц�7D�cs=�������q%�â�(v����^�X7�����b
� x���{�{�;��@7�@�քvw�ηp%�B��C�{7n���>��T/b���;ɳa+Z�i�U�8���ܑ.��̉?Ʋ#а����ѝ��e�M�Ũ�jd�*�ncpc�ޏ��dTzX���A<�u�����	ֳ0+|�:A�ZG^|��.<��IZ��`�t��R΃K�z��B%={���t�V����V��.���N?��w�vb�,7*�K�Ne�#�ie�-������m[��G�u$Nzv���	N5<����=�;��C�Ӓ�V*x��t��a<T��ܻ�V&��:{�L���ՠ<��h�� �6cZJTT�[nK�(�Oݤ��H/�����JEѵ~��

M��x��%{�ad ������cY܈�q�<2FEc�E����3߬�~�u9���b�)������Г6Ζ�'ޓ �D^·��fU�9� L��a�zF>HE���)D(+5���������3p-1Z���o~��{I�&��X|~�a}�p���w��� ��F7�*�����|NCC�ݖ>���s��c��Bg����Z�c��V��:e��e=%�pּ�����Ik����<���}��7�ҥY��V3��֙���y$�[RCy�Kֶ\��B�� i�:�X���
j����[td��v[���D(Ŧ-�10��i�c%�jq��a`�ɮ�B��P�ǐ���(ݕzAɬQ�?a
���F�zl�v������I^3us�#8�h�ޜ-|��%����\n�U�LA�{H �t��̫y0�.�a�E��
��5F[5,�Bg��n��>j\���I7jsYT3a�ɰ�B���U��G%�Gfz�cs�rc�od0��Ί�]la��xQ�+c��LL�af~���H�J�29�ǧ01����+��PSS�Qx�*��p*(�3��%���$ӵ�ђ-^�\~��|z����^���k�X����B��::i�_�# �N.��b�.�X��yE�x�OԮ�o�blr'o,��Ɨɜ�ɂ�-/�+n�S+�8��+�W0���I�q�R��y,�M��������ټ��a�ay)��KE�ͦqs2���Uܚ]���*\�""M�Rf��Ӹv��T74I׋����dyԋ�V0G�k�|�,�|6� �Z�����;�t���\�iB� �B���]䯨��Uu�X!�(�R�"�+�s� ��������J���y��C��$����d=�2鰜͒��(�V�h�w��%�ir�KmҢ��G/��^�#����B�f���_�j��IK;y�0���arfWg��g��T���F	4�,r䭩�4nM�KS���V��&�y�Ed��11��k��ֱ����b��x��$N��DEmQC�'gm�j.�0�r�JCG�MKqK7'0N���tS+�ju�\����
\9��r�KY�O�7����<�[�nZ��e��e;z�;�+S�(�}��g��D)&
X��9����2�[��2J�>�f,��u�08<@�����K�s�@v��~�2d��hY]!�
!�&�	!�K+�zMEf6��
e_�4�Y3�d�~$�����I�����951f�LNߘ��P�Qf	baܿ��=�'�F��|��8�~�j����0������u}�,ꯟ�o��&�Y��ގ��:+��X%�\��V��kJ� n��	K ��{>�#� ����7><���գ>yEaꞃ@<��C�Um6[_=;�~�.ΐ�12Q2������0�ɢ�z�W��ڵ�!p���sp�m�0���@ �������4QT�4J���*����%<���x�os�4���M�fg�e%tӄ�}|h�h8����{(е����&]e�֏�nB80��oC �A囥'p�2%Z�v����'�q� ����5�eL��8ZԸvR�{�k�c�����0�ک����#1�C�W�B%�E��!#l�ߍ_T�==@3�B����NL�v� M�DVSf�hO�k�|�V�R����Jو�F���� ٞ���m�P�Ҡ6-NB=4Ńa?�iK�w�qf+.S������$�n�JTs(��m�kVz�+�&÷�}
�J�$oU^5���>�a��5��]9'-��V)�����,G�ًt�I���J5����+B<�"FA���*�$*���*��N������.Z�j�jG�z������-�jͩ���&�t0�%g],)p���HC-�Yd�7i����BV�y��!F+��|���'��De"K�'D�Nj�@�VZ����<���:���u�V�V)w3?��Y���{��ZNDV�5���L���v7�	Z�Ҷ&m�^"-��/�(N,�
���g�������Ae��(-�:�"y@c���^lHRɰ3����X�V��%���0��=jUDW��b�b�,�lY�,%��GZXO�(@AQ�EUҊ�-Һӈ����B�*ycq�&�I˲VQТ��Y��Έ8Y�K�'�|)�c=6�7����4����
��)���2ή�P�.b{�V0�')b����iZ$��ʏ��z�C���q�ݜf~����C4?-�(����nSR���E�D7�i��E��Lw&;0B ����Z��CZ���ǘ���$���o�ك.֓-�u�T&�F!��Sq���ܲZD� YEE�0�)\մ�Y��m�mN������;��5��V�ڼ`�H̑�����[��_�~3:�^��=��??����Q�h4�O��)|淟ě�u2�&�L6q��|��\e�1??1�#��Z��K�0�o\��M��%�_ɡb�b�) �Q<
l$L�:��-Ody�vX����)��K���-i% kQ�����<�C�E���M{G�,�$��[��߾��K��>CI��^j9��.c���L�<��뫼Ҫf�tL�RG$�_��7a�=���ق.M��򋙵WO�P���������їi�ab�D¬�.,���H&�"� ��j�ꨢ �:��|�Q��px�E$ʊ�jP0i~�D��Ԝf%[eJ���ŗ��gi.v�Y���p�O��D��Ma�p'����ؿk��|��LG�h!�b�A��^e�&�Q�����kI7^�n��;����,�A�w�B6WI��),��G�y�5�Ĵ*\�Fh�n�5�5�̨�MZ|ں[����~4���w�R'X4(�4��&�Rm��Sk�X[�^+WHk�2���+r>e:��>��h����f}ƌ�F��1*����U5��J�k.����6���ӶF&����*:ƥU-��^�<�G^jBa
amgѤ S�T���]UV	n�򗦪�)��y�`��%PQ��)W�7���;_ͶN9ۤ@y5m��|���Ӥf�a��
�)���(���kt��V��<'��z_|h��h.��~j��Q�Ј:�2�|�'�<�A7A
.�Y4���2iܨZ�5��*�ʊ<�x�ŁE��|�t�J�XY�ʂ���{킪�j M�BX�S�a($�$+��_��h��W	�_j���)�f�3���x��	���AZ.�_�G-�m��q��W���s��:��TΠ�'�0�b�&����H�#�d>�j(3��u-h�{�[���(��d2�UR�����*<�<Z��#Z�*@˔J���4
7Β�9D�I��q�:)�:X~�=O�/�O�(.�!**�0���z��<0R*����W���b�_���4^�밗�e�0�a��(���@HL��ן�����X�e��*0��Т�.�2�K�޹��[��@z��W����Id�/�]���^|�?>�G�D��.-Ա�ß�d
��n�����`}X
d�\�����p<G���K3�()��gzS���W�%+*�-�Oc��S,��Z�X�;��Ct�:ú@�Q*��>���}���2����Ïd��%�OO>���,5�����k4�-�@"����II��^lڼC��HuS�3�y�eZ�C�2�4M�)�<vG��4d��4?jk
�Ņ%dҫ� �W\m�Ì�]�J��Ud�Ҧ8�����	�j���XKIS�z^Z�I��i�D��/�0��Ұ�a$Y�(FU
�h������8���.ܽ3�
�|�,&"���'=�����+U�,	�{<y���8ݺ���oa*߁`����o�鬒�e�!�����7�`B���4��,Z�Ϛ`�'߳)%ȵ���&R�j��V"�=b
k��\�iF66�q��*�!	:7r�*��$�=�dnj:z_�I�-�&,DO	��Z���k���(�r.�^E�_0Z�Oۃ�meNa䀠��0��oG��V̭���)Ԍ[a��@@����TH
i.�F?�{f4L��T)���Щ�@�W��0�$iʹVEu@���Ơ��GO �:#pV<�uU��	��	-U��H� �	��7�;^��|�[7���:���)�J ��VwP�{赖���_M��2Jv���d��)��̬���X|����ٖ��B��&g�F�9 �ϕ-ˠ�L�	~��I+W(�y�G�SJ�����$*���o� �Y�>-WE˳�%�x?@K%�;th3*е�#E�͠bȸe1JT�5m�I�d{�Q����Q�6���P{�m�4�&僶KA0J���z�A��"O��d3��2�/�!eŰ�-.fq��̜�:;HF{Ĵ�b<J�a��^�ǋUL'�X)���������d��,�n�._Ň�t^�ƅJs	R	me��G�tV>���#�!?���3�P�0K�4R��;���c���GfJ�+��|����� �]I�S�e��o�ĉ����E������O=`#I��w��8������<���V��{v�͛��U���3�����p>W��!	|��Q���Nu�\��(���?���/YK|(���1g�� z�B��m,���<i#�)�ĿD�����H�Y&��)h��h��%������|�9Z'2���]7�}c���E�������y�6-�x�4�\^�n	b��tz�����~���"��['���"+��O�F��d�+�V�eH϶^½�z�����t�@�fm�v ����{X b��t_|n7'U��,
�toW^	�wm���{���t��/�<��Ity��^�5�ʌ���N
���`/[o@���趇�U�rbѠ���FH�/��Hk
��"�'PPX��dZmf�����%�%��d��i×5�F.A��LL��B^�JBAB�F!P.g��Q��)�I���ۨ�I�����'$(�
j�-j�Z%A�٤ �l������- 	J&j�
��[�ȵ<R�߉^�|���L*��J��
Z{��.
2_cF�s���By�z(���ޖ��=�����P���U�u��˪��t�+8��Tk���f����n)�D#�JBC��j��B��%t���aM�2}�����B��"���B�֒@f�(�.�9�6�#�fZ&j%�3ߪ�3�h1�.+�h�0U���>� UM�g���f=��(����B>����c@k�I�g���U�B��,�L@T�4
���r�Z���`)*~
}��a�����z����}�������r5c�SfrM|�	�Q�SA�0�	R�E��<5���M�I�W��@D}h䓀��%*K�q�Mttv!@����j&>��1\x��ضu�����l.���R���57�E������0��C�b���f�@wf�)d]�K���L�cP��m��U!��ƫ5��#`��k�����<�����x�R!��l{"�Z)Վ�$8�{� ��[v�5[{R1���e߸���*x�&�{w���i�89�����6�����o�Յ�Kk[�1�R�_~���_�Ds�R���
x�n���h	|��=���s,/��c�|Q�N�>���y>~��r��$��mV﯁O�*��~�c/9�C۶u#I��bE�M�c]e	��+�殡�+"CA��K�����AOW�LF �O����Ǐb��lپ{��7ƞ�����G�Y6����,LOڌtY>�H�b���X��Mw�`BY��%��Cf��K����][�p���C�G�42E)�k2&U�Emd\��4��Yn�{b���
N&�,����&����b����O�Ǒ�5t�s��X�tLW��Ng�xu	o�����7��{��Ά^����&�#�c������YB�I��j�%�#���J�x(0����f^M��t}Ґ�9K,Kx�iQk�i�gY"�	�+Α0U�]��� E��e�0�`����j)�he��!+/�IͰ�e����.���8��-�"��3��aТ�pR�������\�&8�,�2M���ʇ�7�O�/��F��d>��`^�Uq4�5K�껊�0e%5ԬC P����N-R[�(|�2luZg�7
�fFz[�ᨩM�"��65�xi�k�� T�n���Y���CbX���	5I��IM^�"v�e��|*n)"��X��*�bC�b�*�h��U@#AeR���\���5eI���b<��NM�$��R��m�,F*Xn
H��N�@�P��&C��� �;��Y}T�d1�H�D<��<���ڌE��F�
��[-P��ڡ��j�Y�T�+�T�r7U'U~!�-I�+m{_(�����RV�����DH��^�U҉U_���I��OZ�h��(?l�qʆ +h$6��C�q��U��c�h��Ӌ��<�n�#3�F���Bp�:{q�V@�K~�5%�fm"Z���H��P�z1��E�"�ky*�u�����~�1�j~cy���M��iî�1�NS��G*�8�N�|�m%m��^�����=����	��3M�+�'=�r"Pj0�u|����G/����/�� T�|��r	�:r��U\<�eT��Z���uն�2��o;^�w�Ϊ	���Z�cײ��WlO�9�%pQV�5��b�S~�X?��	>� yV�L��g�S(-R�(`j̠�]G��M��OG=�J�
��W1GƊ�Լ��y�60 s�4������Wp��)���bhx=�����Μ>��g�cii�[^G,�H% �^X���i6Q1��o��6e�g��"Q�<��K�k��>��݈t�!�9�.f0EbМ'��[~�K�O�4�S��cV���� �^Z�zw4�=[�(d���p�2��[��V\� ��6V�X_��������q�B�Vp��go:�(���(R�+��L:-�Y�u�����?ԯ!M2Ҝ$i�j'XTlyu����̕b%/���k�'�JsT���i�Li�T�H6i�-f�К�P��@�0�s��C��`���⴬"|�t�)I#�Ĩ5j9��Aq��RӐ������.��YJnj�N��&�|1�j�QqJ��YN�;�&��P �x�Y
p�Lֈ4r���`b�J������	5YP��WUs	k���qKp�jSв����W�U��,2�ɏ |����W�꯱�
]�?M\�[���T�j�X�j^r3�N� Oit,#��<1QZ�^�G��~5����� �k�$��'`�E�Zj��F,o�ʬ۹h�,�K/�`Y�(P��>-�\y�u��� ��FJ�j��o�~7��L2_�W��@Re�4��Y�2Y�	�O���7���J��j�14K�p�d	�iˊTZ4���Tv�4ZR⊋|�i��Vy��F *��y~�s�2߲�ȇA���m0�J�de�l�n�a��14��T/�����a�eJ������ ��,�o�e*Β���2�3�~�����VJn���DheP*+��J1�VI�eu2�2%�ꭄ�õ�E��іwmg�*�7��VɅ����mí�5�M�v�C�W�bxח
��g��±���TX\X�T�ɗn�o�t玬0LFf�jA�1"�#�`�L�s0�:f�Q��
2�%�[SV6�6�P��l2����t���G/���!?{~�������(�Y ��I}�X�FP� �e�]��KX�ycY̭�Tͦ�ϕLs*k�E���K�3Ճm۷ch�:����`2�<�$�lڄ��AҴ��I��>���Sb8҄ךd>%�=�j�!/�q�:�����k�|;܍ѭ;�~t�׏�whɾĻ�I �я�7nZ��uX��"�'C�����[}-�ػ�Q��<���	>��1^OC�3j�
����L[4�����0N펐/}��C{�S�x�ٱ� �V�P���B���KF�~
a	�5TM�ը�05� � �ײC	/Yr�w�f
�0'���	t+q	^Vr	E13���*�MM#�2��2`Z�\��Ț:�d��:5�6)T�s&dZL[���b��e@ݖ �Qc��]�i��A��-@�j���z��%��:iaA/� `��f�vc���3_�u��A��jR��H4���ey(<7�VyiUu�Q�i45�A��Dm�Ξ��3s�[J�UM�Z��@J�#)e�����u+<Y��gSe��-mT�{^�(��X��)ut�4�����g�A��F��i�J��C��0�8�����\i9-{����R�2Z�K`��4������+�2i��.3�RZO��@!],�J��,��6(:��8H�7��Ls�h�r�neuSHљ��xV��h��)K��<*-�Y����4*��a����F�9q
�.V?��5�X+���/�4A��J�ٶ�,��%]��0��N���K�2I�`r��^h�B�R!�(�!>tk�p	|�g��D���Y��*+��NW07QG~��D_�T��&��y���@�i�S�yI���� �$*+�u Sm!_a��Hؚ�ֱ}.��Q��k�x^��D#FB�3z1��Ъ�=��n�\�t��.���*�M-Sު��h}��B~�_���b�y�:��//�~���U*�ӬG�;;��|�2��H��%x�(���H
E��w0���,It�S���e����(WP�|c�;�[H�|�&���RM����c}�h{�@2��2~Z�"�Y�/͠z�k6gB����e�Fl�8��u�رc�e�E�1f2G<��L�_#�x\�d�^^Ʊ�^�>�w&�4#��N6��V@qL�3B�H��fEMFj�u޹k�V��O��;���rV(D�MA�>�J!Zc�i� 7&����qܼ~12���r+�FT!�)�[	l���>�w�فy
��?}	Oo"����a/�vW#��l��2l����]�{���x�Hu�X0V�l~���H�
�z��%ZE�F��H:�]�i�՚��U�%��m��U�1_��%����aİ$dj�'P	�D91��2(�h]Qxi� @<�Nm�/iwJ����P��e蹚DC���1���kͼh+��D��M�B"�D$F-�����j~�
xȀ�>ԏ*!��&Չ�QM�8++���i��/�Vc���y����B��1�f�CeG`(e���
wUv}g�>̋i�̛�!
��U:=|W��e���>���JC���rd�լ�!�Gۀ���:����:�U���h��N5j�̸���aI+t3*�~*a��8���9֍E��V��Q%��&�ު2�򲬚 ~���R~��ZD�S#�ɢ
[���Y'iQ͖��W��35-�i\�,P��(� �[a��<A����A�:#�1$�`����"���u�{�YM� ��t�4T�i�3(�H�%j�Z����E�]���/��V�e�Q��\�pr��H��� >�͚c��N�R"ͩ���Y���Gj��D�(�"�y#�k_���@�1?���A-B'1F y����e���i�Gh� On���L����"[��˓n�����7��
Q<��8k������	�H.��FV�&��s�JGY�g�&����s��X����6����eD^͸����^9���g�o�2I����k���3�+y�E��� �8H㴴[��'�� gu�갔3��ʂ�����!Za]���N��U���� ˋ_�C�V�H�`\E���|���sI�ݘ�_��H>��4Y#�)lmeP:�4.M�b�N�TkNql�0���v@��$=��C,�ht��'/������~��#�Ȕjn�0Ғb^����\d�?+����iq9����ï{��Z�FZp��%GD�f��4����,~�w�Ǐ�B+��	+�oյ����J9���~ܷ�ϝ��o���K-���0��!jo{�bt�6���:Ӵ�bHF�ge�Zf��5
�B�bj�%�l)��E��]�5B��4��+_H[�ج�$��(+"5H	���)&�ѴOsu�������E0	I��)l�ɗHwY%�KMr~�O� 6A�
bV�J �{Һ�R.�1�@����Ny��(^�Je��*,1_ �t3,Jf{ �Y֐�@��J U'|��Y�>����� ;::�81��O��u5
�F�1��#	v�D��OM�j/�5S��QL�v��6jr*�3ˊ&0��Z�s�Q�]������b�
��c��B�G�W}r��X׀
j5e�yn�����G��+�V�Gjх*ҫ��i��,�)����9��LAԶ,�"�J�/v�:�o�(�+�+*֚ ˬFb3L��>.5���piر��<��)�#k�L���EL���|�^�C� 
1R��WZ,yѶ�W5��������N�In
M5��g$v����U�?���6��VNv��idn���E��G�U4��zB`����g�^�"(eV�6��|�m3B�8قJ�G��+Յ*�H���E�:[�H��-ύcj�nMO���[x�L�1��i\$n+���=BE+I�2@�ýĄ>������*%�m�!S�(a���,tn�@S*���<��6��)�?��ㅋr��-�Wju�7e��*�a�V��;ڥ���,��1���x�MC��LkS���za�����8}n.Ҋ�Pmp���x�T�:Z�u각A�����}><�h��R�e�� ����>JB��´p�"���j���Ud-��F�}�,_]��L�&M�I$�on�+x�/	L����"A��J�g���p��؜�-ͣ�s ��� �p�
5(F-S��Z���]a��������+X�����I9� �B�38�%��#�
w�ڈ�����׿�h'+;�^VZ?Y�,,e1)&�8�5\�:�O}�s�v��Y�fk$T3�0r���غ��y�]�k�N,�����F��}�I��'RxS�(�r�6&�����J�t��'m͒���<2d>.4��A�����,5<U�:�k���,D���WWQ(�,�e����
��T�54��1�:�ɋ�� [����J���,U|		41�ĸ��վ[��b�G�t(0�,��(�HcS?�x�J�RM~Z���I��*����6G�&! .$_�G��h��yN�t�7�UZf
�L�*j�V�,5�)�d��̲�)�BF��eV��	Q��S�r�<I�O*|c�}�J����YF|W�*i�ڕU�����"P�Q���yA�
��mլ#�z	�xQ��8�djMi&aG``Yh��@9���~ӦQ;����V��~0�L.�r��X�%��-�P��JQc���&S���B*��d��gU���v�Qc����n�Y7�"K�����h��
ѢSߐ��ڴy#��@gqn�p;�XzW2e,��Yo�P�� �w�6O�_��Rc^eA��0UH_Y��ڛK���ʴ&Y�3i֑�\�"a/i������e,�G��:C%��4��g�(��.�=���H6��>�a��Jtm�?�M�1��*���.��Nl�~��ʭa
�3/���/�G_�3Uj��--2E���I~!�EWh5�H���!\M'qvޏtE��@�/���ޮ�+-*�f�H��3	�6�HQ�\dYJ҉pRn��X�Ь���%�]Z9jr�Τ�,���+�}�b�1���;�q������F$B%�e�����/O����7�^�ҩ%LXwe�X��d�ȉ��%*Ydtf����xw��,g�j�AG#5�ԡ����/�\�!�b^(��~~
��=��k��	>.�P���x˺���a%"�ZH#��!��ʯ�k�g%TEW��u�E"4$�XZ�Zp92s��T1����2?-,��֭I�>u
�?�M<���)�w8�T��$ם����܋7��Q���Ѵ��l��E�_Z�`!�J��-����o����Yj�ԀE��T�қ  �u&��&��_s w�ݍ9
Ǐ�r�^8�Jo
���^�wm�}��N~�4�*ר]�\�(�V�}�O�va��\�Y!M
&,,<mP�6T5��rP�y�V����
b��~�0��CR���bni�%=U�Z�����Z�&ZB�/�[Ҟ��|i5P�O4�S9�$T1�	f����#<��	�zQ�=]� %x,���H�&�ժs
&Ǌ�Η�n��+���g��"�j�]N����j��:�;�:)(i���j*�̃3�Uj���OxOWeY�Pi�':	\�fi����Z�0O����&'5��o3C�lÇY8 1�0Ԩ?�_�,��%�� X�%/��,!�eZH�����6�D!몫��o�֛�ayy����C돖�Ff��x���d���:�݃UN!Z�]�ݖ7gd`��dm�M���Rpi�D�uO@�z�fX��	RS�nj�J��f�T�������4�P�kT�����&S�	Fe�j�)C6\����Ӱk��~u��U�F���mM�V~�OΥ~�-���d�J˴P�p��1{�:Z�G���ʲX_]C�e��@d�L�Gt�a{�K� L Z%��/�i����?�m;6�#6@��ܙ��=_×_9���KPt�zj�#T>��^�����pX/�)�=��.���r�FJ^3�u�C/��y�i~s�m�i@�g6���Iaַ���)~���jD?�VV�:�f�h�;��6���a�r�T ͮ ��}�^��P6tS}g������w-*:���ׁq�`��S�#f��U�*�G�ki ��#��Z���d�
����M2�5��D�|��0�G��|��~�ϟƒ,/���Q�ؠ��R������E�2����$ɨ�|�HiX$�� �� y�>	U�\6o���Q���Oh�H-�ި�y���"�n��_�{�՟��1�N��d{����R8�w�l��5<X�R�:�(SE1@�)bfv	�N]ƍ�& �����N7iQh4MA-��e�?�ڻq�=�`����I�=��@ɮ>�a/޾~+�}j�H̤4�Rc;����'m��I`�i�kt�4G�%�XJ�
�3j�fq�#nB���eŨ�-�#�z�_3P� $8��J� �\!
�����@�g���Us� H�X��c}��(�*	r�	�%���MV�&�VJE2[�B<��M��(���ת�	B�*/�e��tK�S�1�P�c�d�D���zVY��G -���,K���4Ej���%-Y�%S�x��x�u��5L�*+�{b�[���P�DLYvF�O��X���	ֲ5�C�+%J��&Y;��эe�Z���<X��t��'�?c��J��M�2=>D�w���&2���٣��
�N�'�񈄷�N�FJY`^���4f�G) �.��7vT�̿�[ui��)"jH��LtR�4x� �!"���u-��Q��wt����ꭽ�s��v]n{��y켷v[�$ySM�zH���+�R�&��cyfS׾��cgP^�"od�Z�bA7)Ҡ�V @�]�=��Һ�Y_�YZ>Z�i5��؅m;���w=��E\<�<���W��S��l����w�EYaYm�40J[�G+��Z�M���F?.�D1�S�	�������".�D������v�s�*��
��ʐ4U���6SY'aȧ)ҧL�0��|<y�W�Kuy��u�x�;w��ވ�757�_^[�/�{�����q������cf%�6��qD~�d��y=P���z��RhR��D��6����ފN��o�Sgd�|\�g��������.����b�j�V������� |$��z6 Ą�yG���В
��M@)R�2��Z��i�RKk�R+R�0���X����
�����~�?�ġ>T�%8�W�Ja�
@ό[�ċX=�85Y	2K��e�%p4�nu��ٹe( ;:b�&�����	3ci�"ض����=�g�.L����/���h�e�߿��߀�;��F�/2�iV�`��idX)4�B�Ȥ�#߫���3Y��`Ĕ*Y#A
Vm�ܑJ!O��3x+��kN�~�9Dp�्0�6��NE�d �zW�0,���H/��-��گ�,�ĭ>%)a�4*#}`a�#�����~�����V{���g��w��"T�-=^��5��}��R��P
Cys��>tB����"O��7���{5>�LTY{fD��^�wGtt��Uǵ�r��+��Z����ZP�K�����Ļ�x����������*ݔ��&�9����r�ǹ�g���Fg��y�޳���N:��۴shy۵	c�o�����5����D�vk�S�RiY�VtM,R�V=�r�E̍�J�B�*�����}�\c�pSĻ6Q�OiG"��dJ��:�ؿ�(�q��3x��g���'�l�u7N�;9L�'m˾�ೱ�Cty��S�Io��n\LG���}M�7!��<�'m����X=m�i��')Rd�������A�My�3�^@[U*;�����hI�4�C|�����=��ۊ�b�ʠ�OM�Kg��Q��&eܘ�bl*�.M4i}��w��F�3gNVT
����t�o,Jջ:�Z��i��0��Xx�^�Ff�|	 >5*T�����Ї/O��S(.2 �/K�%0�J`�FM� �yBӴ�D;�3�ry���jqy%MM\���2ZMe�Fh�K�T*4����/����Y���=�_��c/�d�w��_e�����9�I=�e]�Ůd�_�`n>�ZRS���Y���Agњ1��o��"P2�֑�t�yh�!���N�7���@?�L�L�N�����n�%��`}��c�g�Hl	���S(�	�b���ТP�V�v#�9�ޡ���EO�FtlD���nE�s=���Vz��)�d�l|�,Qzq�Q���2k�W��[���Y��q�ѵs.Z��9���-�ݵ#��5��Մ�& �)OA����v�v�pפb�;G@�q-o��~�k>s*�^ԿC��[��tw��s^�r�w^��.���}�A�6�� �|;����V����^e N�t�9w.%u����ް�$�]���8[�Ў�p�����3��g��#K���9�3{C?<8���V[9��Nn���:�k���^���5��r�����Է`�̹	Eѷn������6���!�L"���dj��fu(S>d���/�Q�R�)�b��I���^���9ZScS�>=��%�H�0�&����$*��8[ �G�p�P��\�!��[2,��1:)Q��+v�r�E�|�IhM�:��{�P����/���yG�b7N�5̣V���:}X�� ���=�������٩#]hᳯ���,����_���x�cUk�O��f�v�K��R㋶aw,<Ȣ���R���G� ʛ6�*l���\����Pm܂o�1�i�(`
�t��b��@wѴ��ڣ@�l�V�*�%���������ZI�`��[�q���x+�k̕f�AS���	PehD�u�2n'��m�+�f���^
d&��U	ZDm��1��A�*�|�r��
�������#��F�6�N�g\���W��c��4bJ�DA�������2��e�+4�5�J�BqS�gzl�2�і���Ҋ	�{��݈���08r �C��߿�=�ll�.k�t��ܐ������N�'m��;��^e&�1�}$�г�:4�c�%T4ҳ5S��Vi��3^hb^�9qhЀ��;r
ɴ%Y_<:!;q9�nG�+שnf���[ʇ���?p�sz�s�g�޾S�
����=[f�b���k�:���N����}e���v�i���󖽮�Oik����b;(�t:����N�*9���y�i�dAX=���%�(ܵ��!�=u�|�_������L� ���=s��������{vq�s�ඳ�t-k���g����N9��c��<�������a��;��Q<�rl2԰��0Ҵ��sW�;��� �J�����kS2��(�./3��=U�V�|�@#+m��Ej�>4�Rs��̴��g���_%Z��t���f���u��kk5k�;���e�+0L-���Ļߴ?����������񾟹���{�?��������)��@�V]x��4�䣧p����p���C��!cIe���;xZuI2\�pʸ�xCWk�\�}�]eYa�'8+b�(O�u�X�:�]�y�N۞L+)���m��p�f��bu�y�W�:������j���Hs7t�A+]�R,D�\1O-��NMv$�E��BBP���D�Δ9ް��.��E D�h�3X�3[�� ��x��A���fw7<���H�"�م��~��t��dZ�ͤ�A� S�:���ϋ
�U#C���H&#�s�����E�	>"���8FE���i�k��F��"�܋��bt�!�p��n�E�/by�)�Ѥ,�\�ѿ�u������S��m�k�pMp8BA�������&̇���p-��{���Q��uR��G��;?�sB�ӧd��I��o���?�s�8���ߚsΜo��{́p�8Ι�a*���ZHv4Z�����v�n�}�'��=�����饸�y;�:���vktp�]圼�E�;��	�W��*��u%�b�}z���N�,������gu��2�G���N��s���=һ�w����vk�|����㑕���n�q�Q�׊����B4��#>�׽��Dסآ�[Wr/��=(����F��
r�3��'\¬�Rx�M�<"���&�Yƽ�8�e�.k7A�^S/	!���J�R|պcW�ү4�GёX����@G��=壛iq������b�����/�w?������n�o�}����ߎ�����ۍ��)N�\����z�,N�0Ƽ1��nz%g%�iQ��ZZێ��v%N3�4^a�x���p���\���w_u���K���3_g=Ò�q:�2��x�H�n9#��l���%��Zؚ����t:�`ZHt���2-f\�4jI3�"j��3ឈ�lD��eǉ��d��Z��L:��>�h����ExO#�H���?0��L_-�8RI?R	��4ڏͣC��LZ�T3��)m+-�kh������I��{͑Ђ����v.e���Q/�(���Jy�޴+k�{=h���ۇDr=AY�q�a��7m�d���G�ǎ�V�w���B�g���������:u�u�	��?��Ĳ�n���������g�M��Ͷ翡�s.�НI/�r'���qӿZn;�J	]{n����"����S�k��}k�}g���������C��v�����gk�}��H3���v�4�ݕwZ"t_�V��L~�{�O����j�r��(*N�ng^�IC�a�����8�k׷�����҉N���o2�����&P�^����"\�x��k���n1��?�-�z�'���{�����V���p����Pn��K�X�,`��Oֶ4!][�t4����i�Hj��J.�M�)���(�֧-9�&s�2u�x}g���hu�<I�g�Ґťu��k���~H����j*�j�+�71�b]ԋ��]n�F4�Z���I�e��5�i�`���Zdjv�
_�\+��v�^8V��ٯ��;�][��-o��K��ū�c��+�h{	-!`Lŏ��v:�YHjF�e�p~K`q��:���KG?��l&�
-$u�k�0HYJ`r�t�~<B�/ALBhݡpXC/}�$�v�̫,mO)��a��;@���?D�!hE��U32�Kp�ņ�I�P�At�0�b�7�-�z02؃��m�k$���!�d�E���if��,���J����0kP��˘�.؄G��:�ƴ1�-W��v�@G�6xB��b/���Es'ok���x�*�Wo����M]�{���n�_�[�T���Bwb����N�gm�f0��c�	D^����N -�0�����{v�0\k�9��s�k�;ޡ�ܫﯽ���B��q}�[R�|m�W�q��m�kܦ������զ�yi�w��;�A�}+E�	O"E�� W@���j�V�����r��r����[�[P�ч탤B;�k�-.�޹g��GWk�NK��U�(�$y��6G;n-!t
W�z�����k&���Q�|Ϭ	X���i���=��q�#(�|�S'P����޸�۶"�RS{��?�3�W�V���:ܝ5��8�5���NZ,�����5Y�I�$c����N��)�W��&oK0��V��\M�I�Z%�)KJV�Z�I��Z*71�X�ߝ�����e|���t�*�}��\�Ʒ����8N\[��r���q������x������-�K�V�2�&�I�6�Gw�v�up��%ϋ5O��|�9ŧ����;�����Jܹ����ў���O�Dq9���n�-	�>8ԁ��IH+�C������wi��#n�n��1ّ����h}2EMhwS�[ZAe
�j�-�����'O��S��ɒS1�)��7�	<d2�-��sM�}HD���4�AJ���Vȯ�G�y������"
�*h�����F@�Ū���e(�ޞ���NL`&;�V�D�eȈ<:��� ��CU�*��x�]��D�l���l�w;/�dk����NtZ��k;#S�pl�ԡ�*�8M�W災o?m��w�����)�J�Q�}�*U`G�ur��vl�����F#^�QXN�n��i2�KN���?���4����UOo� f}*^��@1�Ezy��71y�
&Ʈbin
��sȦ��i�k���T�NkO���+�����j֟��S
r�FJ{;��*�D�疰�0k}�ɮ��I*�uԫ��6ܵ��D��*���؍[��Kc�UAU�����<����tPy��Q�3�Dӛ�jم����,'�\)�og_��=L��ӱ<��-����FoI�ڵ�0W�40�)��l�n��+�x���??��NL���`v5�$�`g�2�ud A�2��7JU�z(�S��)����4�I��I_�JE;%�ߵ��L��M�TYkZA�³^7=km���C �s}n�Ĭ@��%}K�ا�M���i,]^09��G.Z#�0#���o��͏����!�b��:۲��i#b���<5wh�41L4�6?�%F4ZiW������2斗��q}�&��կ���,)��2ݲ��LoZ�NBJ+	�`A�C�P^�Ei3+��d�z�58���i�*B4w�Z0MV��S��A�g��Jyjm;O�$�cx�#�q஍h�����s86�"j��cei�7�z~��?�`��R�*h���# ŭ*�ל6y�G}=N��o�O;	\�d�nbtq6�H�O���QU�dj	\��ֿ}ga���8S���;�F�k����Z�?JբmM�27��[S�����'H�{����3��62t�7��<,k�j�������9�ά:ɟ;�4��:U�j!X����Kp���8sy��Z�����P��b�ژP�BJa8�v���w�� ��o�z, j�<<�4�� O;-�TX%�P����ٱ[����%DU��s7�!/j+PZ�
�l��ѷ�t�4e���Sx��#x���/f0�+����@(�(󶎊roiqj���(r�Ǖ�:�ͺ�P�2�j�S�W:��I��Y��h�	�z�e�����I��$���WSVQ��g��$�2�.���yq��ZXR]Eާ�mR�!E���[�^��F�l��U��ٙ�ue��M�*._Y�S�_"]i��p(�&�T���j�xlXݓ��|G8kx�R�a�����=�^~��6χ�2�P :��:�V8�->���\���n��Rt��x��xH�&��a�<�'M�"�j:G�E�6��.� ��2'a�L�f\+6�����X�̧	}�l�l�s��Z*Vp��ǅ����
��P�uf�F�pU@�^�K�ζ� H&�
����4q�P�Qq�	DV�\݅UZ:+�x���r����Zn�K-��Q"e�>lN���5�[�+�*�B#\`�r�ҍ�����m���-]ʑ�@3�vV��d���_^)'����v���S��H"��h�)um�S���I�6���K�����^���N��5��)�ox��w�x2�<.�}/<�5|������~�z�9���	���<�܋8z�(Gm��zn�	�?U����2����m�i��Z�&y�� :������ѿ�>�������&^|�4.]���?_�&Pkq�b���9�r�Μ��Kg��ԥ�x��+�x��p�V�l%	��MSv����?	r%��ڣ��c�x�̭��HR�جd�r���P�"O!���T33����D�\G �@I+m�R����X��-���2�Ez�yo.�DV��$�D�;h(j�ӥ	�Z-B�)k�CK�W/�@[�ޔ'�8�%�Byl�ӆ�3�R����j7ف4lVY���Pj�SE�Tk����"B��a�P�t��h�D_�p��� ��������`�NEc���J��~��U�T�[T�]T*�Hi�;�-,��̫���2�&�k�_�Ї>|c>�ϟ#�F�z�A��������ؓ�1�+�9,-�Ь�7�В\��I��h�i�D���?`Kv�����f���`�Z�-�N@�����
�:n\��$T1��B-�֏F���ͭN>Y=" K�$ey�#���}r��2��+�5�$�e�+�I����:�Wӄ4�V�VRW[F�08��{^\_]�Tn��yPEs�ډ{��!��s�ـ�Ť�jm�Iy3�T:�Pu��։Bk��AfU�4�z)�ى1\�~��C�"��_����Um����	���n-�m
ع�4�K��⋟�4������:���p��,F�ad�nt���`|z����q��e�>q+3��v!� X�-l)_�y�����6z�7EO�<t�V�.�?�?��?�G������}/9�p�=�&��]�Ż��]x׻ގ7��x��O�5O<���?��x�ׯy�B�V�מ�N�>�SW���/A����p?��.�iòը*��v�U������h{R:}�Lk����c��:C��h�~��6 �هZͅ��i,�O�Q���p��Y��2D�॥���-���u0ҍ�'�t������z/�$��N��=L��e�Zyj�jj}�B��-x�<2}.Zd-����CRY��� )�4�S'�BqP�i"�&�JȻ+xk^dsL�k�Q\źx}]1�I�A&����|��e��
��[�J'Ot�{�㎼�̚�g䶤�xNyפQa������4��C�}s��la�n��e�-_?7��s��D��/h��M�0Q���w��xp0E�g�H1�w��ݽ�d��~�2�5y���"Juh��M4����*�iu�����#��j%rLL��o~���7�J'��&~6C�V�(�$����0����SU��}�|o��L�a� i�������5��W~��hQ!��4)�k3N�(��	���ܳs3��P>u�$�μ�Jr�ϧ1�/�~?��w��q?SJ��ڤ��Rs� K�b<9i�T�|SO�������FxQqXY^�����{\ɮ"A+�o�fD�qtD�ݵ;�@��0��8s���9��ڭY9��������L��ɓ����}ܸy����Cb���X?�]����3J.Ԩ��&�	gp��q<���a�׍���o{�?�6���ZW��R�H$y�2�wNE"+ԑK-��L���O}ߠ���3��ǃ�<���{w���-��كhD��)����ӥ�j��"f���/�����O����v���m������ �I�%V(�5�����3&P�C^a��s�����PZ9����S�h���+~tm>��-�)Æ�)�q���x�E�]:�+��0�*eT�O�p�$��s�az�C�_�#(�⸱���%?*|�Ep��Nr=����R)�x�Z`�i�V���|$v�ٌJ�u�5��RL���(	�?�P��PIduh�hw���C�{\��l���xn5=6\���x��8~����L3ny��yN�-�����9WW����\KJ�2Hjv[^��E+�@���@Rl,^^+{M.�3_��jy�V�kg��s�>!��c���f���j��U$G��mh�w�@G2���UZ;9�����Z��(��'#�0�^[1X\��9uR1�r!���2Ʈ���g��,b~f�����C2�IK$�,	;7�uƅǩ��H�~��R����C�#&`2��"����1��;�k���,\���
 2Kc����7��=��a^��qd�e�:f��8�mǏ�| �}Û�?��du���j2�fՕ�N�нv�~������v��ŋ���|/>�4�i�y�[�o�vtC�.̎ayi�xO<��ڷ��2��Ba����|��[����}���q��	�>ZO�'���'��F��\  ˟�%>'PW+.֙�\���~�[xᅧp��صqoz�[�#��O�o� D�5�7�o��	��M�8v�e|������u,����׿o|�;x֍�C,B�Ǻ�E3����̧��lxF��4���_�����1�y1��C��Ə����}�-W�4E1Em����9	�A�ӟ����/`�]c�3N�sC�c`�>��D�|�f�q��y���q�z�4.P���>7�d�t�f��EtW��vږ
�:n-�0Y��j+�8���K|�SgP�(5}��ծ�Zq2�!ZѼ�������>�@*�W� ˂�Hp30�;e�h��f�����ڹ&�r�7��p�#]�,U+P��R��
�l7&����U(<�F�����ǡ�E$z*H����碹�v�mGh����v�`VX�'�!�L ۇN�����'D�)U[-m����,�o|�@w�/Ě��em��pv��_F�Zf4#�h�l����r�2[j���D�L椚��5h���$AZ#�B�$���8K�z�B<���w���ﳑfWi�Z,�� Z1Ӭl��	�$ʪi�ڄ�ǣ �di�8ϥ=�Q�SA�ё�m�ib���M��@k[w�pۿ˥*~�[O㹉Q���;K8�܊�������ﺟ���',VV6U�#^t��x���F��J���=]������L|�;��o(\%���]�=z�kt���?��9��^V��|xT��Q;,��g���nG{`y���G�Ρ��QH���?9������>����ྻp���}�t����Ղ�%�ݘ���Ǩ�񶷽w�7�� J�ծX�Վ�k��(V����>�_����ظ�Y]~�C����?�DHMQ�yq���:oy�DaN%o�ũ������t��}�}~���G�_�mb(������@�꬝j�,�~�[��?�c���Q����]o{����b�֭)X���!F��ȟ@k��K�K)Ŋ_%ĺ~�:<�"�35A������>�o=�>E�����_����C�_ہ�A�p:��aW�u?}������[��w �p���ų�b�`�q���Sx��gq�[�8lb���&�nZa�(GFh!%�y�(/��V��xJQ̡�Vl�˷�?�<[�;��d��Jx��}�Vz�[���[���A�߃��5*�ZeZ}�aFeY4d"�Y8j�	��g��qj<J^����G��
�!}\J8-[]A�Y�u� ���F0(�O��ȳސ�<����4Z>��O� �le .�
���I�ʅi���,������_�[�WN���)3!� �m�fZ��A�EШ�h*VQ����3�EF6=;���Yj����_��b�X\^����r+4��0�����,��zaK�fqq	镴�)��P��ދ���hUhE߉�9�T��ѐ�&��R8~[A@ϵ��1� �^}?Fv_�N!&��G�LB��#0�髌]��G��q�8�����Wq��M�Z���o��^Bw3�}��y�;6���Nǡ��(g��Ν뵃�M<k�pF�X
�G}��#�ҋ�xmR���~xˀ��#3���p
K֩�t;BN18�v-ls�8�keA�kw�<�BO,�Ι�썵��)�fp���I��=����w�ރ7��ͨPQ8�%��iLMM���ȓ�6cp�(�j�c���k��;�g����L9c?~��o�)�G�G�ܵ}[wnGg��b�R�i��m).�pS��.����G7c9WƱcGX���va�=�N�t��ڴ��2����׈�W�ş�ٟ�[O?�����~����w}֏�PYw�nm�&���Q�K�c|����vY+���q��/�
��9����#�D"���-��g�^D���ͯ<���������w��lX���pTNX���J�J܉��A]��x�VG}�zբ��JS�hP.�Ʊ4+���?
t�ԯ�F����� �HG���B�h2�������J�(/�$��d��N�S}oJ�RW��J�W�35��q�ha�5�M@ K���s��	ND3�1�
T��S�<��6���!�i���s��u�Ak���A
:WX*"���n�kECo(g��]�'엷M�������f�1�Z���ų��>m�u���eB/YfX�B.���n���	�� \�g�o�7;�ߍ�ލ�&`�J�4�hL��کЯs.��c4Na�zSx�[�k��T�6��Fp+�Z~�N�V�:���^
���*4y�f:qE �%��\SAl�r���N�<Sb,�J��0�Xg/٬ٔ��Z�F� �s�<֪��bS'S
�v���!MM#�G�+r2�*���ki�*]H��F�T\�VyS~L{u��;c��^��҉�xJ�:��%�8�>ι�[��󥂲�����)�Ly�+x�ŗme�7��ؾs����$:�~6��k��WΏa��Uc۞�H�r��ڱ�`�����&}�WW����4.]��~BG~і���W�O~
�.�A�Z k�E,敥Gڒ��3/T�b�/{wm����O����>ܘ]dO����s����q�����>�<�̳غ����~O>�z��vS�9���Zt8�[d�q&g[���b}�ƋZi9�����3O=�S��bu^0�2Вڼq?���O��O���1���,��y���I�JHڿ��-�C�;�4��|�"�	W� 7K0��P�o@*j���`�nԃGvt�ёa��DR �-ZQ��n��i�7����l�Ef���c����G��z.G�H|h9�L���l�z��NW�������.*���球?���B"*�kE<xݞ|�]{��݃��O9#�MZ�·(/$���S��z�~����2�H'�Z��޹���y���p�����9i!#��j\ ��y��c��*�u@Mh̤���wý�^�~�0���������oy#v��mıi�;�i�v#�z��SM$��A
'i�����h"	���F�����.�?���˴�|�ڠJ����iਙ�)�������|� $"���u�TN-�)�&xYqX��Bμ4�:-/���ۄ��ѝ�czḅ2�ba<��4���mp�\L�PLt(,VJ��;j�56'�it��S�	@��W�kU΀�s[�3�M���A2K��>�
#1�����r�m?i�\iB��9Ͷ���r�[\���g�{�v�;�D��qy�9؇�{v`�ޝܲ	�T/��c`d=�� �oM���p�M�D;����8G�����1���o��ӕ�9"7&f�������o~���r�j�2y�Ez��ȱ�li(+'�ւ�{�n��ſ��C���+��G>�t{�`��?tw�kuu���g���|��K�����k�x��sʊ��
YY]��_�������{��_��O�l���"��5�6~�����ӟ���lB�wk\D~���7]=x�� x���g���5%Ŭ򲥴-$5�J�H�\�h'�ȌeP[)�UȒ���n��@^o�P�- ���vl�}���-�asl�䢔�zC��:]�(���!�*��%����q̇�Ê��O�z�R�֡�����&��Yz})���ͳ�)<~g�T�訊"�E t8w�Ж$�E��+��I^0@5����W<<�[�u������C���a&����`�������z��v���~���o��J�:�XQ�h�z���
���@�hI��G��k�v<x�v�?���ط#�w�.�N,"F���A��]�}Hv"���k���B$z7����C����N�8���N"�4g#�>�#��~"�	T���įŧK��uC�пԘ��%�6�Ԟ��}SK�Pñ�W�ȗ�Hg�XaE�Q��2N��`w�Ł��H%��t\sNa)N��?pJ� O��
h��|3����,������U�����'+d��6�� �aT�QM��1�?�@����eY�@'�WX�v%"���s�T��7�JѾ�����-j�����p�F6�G�:�����<��sx��o���}�N�+P����A��w��Ba����F�w�]�TߔʕLO}�똘"��-o}+�۰m�v{.axql������������!{��.��������γ<��$볾b��}!�ݹ��!��}��9\�Χ�'��p��tg�iQ3��a���?������r^0f�g������7~�q��et��C���W>�|�s���B������4���W�]G���� �5ӬV�����w�� ����b���_��o�PX��Q�F�'���Ja�Ra��I��Fa���V؟�Qf�p���R#�Gz@	�vwcS_�Stjks
n��,�l��֤�
TTG�[��>��z�or����0URy�$�&oIɷp(om��Z}�=�Zx��������>1@ij�iST��u��RW�L��G�Z^~��Z��8���Lxn+ ��Ӓ��u}�r�w'���68J�Wx���f�Z��<�L�C�LiMO�$��舆ъF�e�0�މ��6��'���8�oY���( z�ё������ӓ��`?�<�B8��!HM��ۅ�p�7a�*@i���)��_B�,ZM��]`4�BM�T�1�Mڰ�*��J�&55?mLa��Z��:}���[�j�}U���}:��2�"��������E�L.`af�r�L>�d3��]�® ɧY�Q�R�$-�8�,j��g��K˴���E���E������.�W���G�#���ק�����:���o�].��C���`�2��������unZv�ʁ�g��:���D@>��\��JQm�x%�Ny��1r�����X>Ñ��L ^fz���:a5�Po]��ų�p��y�|�e�Ǣ�[ᥦ�m�#�+J�:�ۂV%�3w�}n�j�51���8˝��<����}8x�^��=x����_��/�ozrM�8w�����~��q���1;=��W����2;F�Yf(N�%ߺQ<��#8��CH�Wq���%��,7G���6	l��091iS'�?�Z������y|�~����?���������}?���4�+_����*����RT����O
��ro{������O�����>7���2P�U�½��'ڍ/�;��k7(d)�n|��+�m�lr/ ��Zi���V)S��*ʔiM�rܚ�˴>f�s�v�.��&O �ZD%����f�7�P�SJn:n�^k�r|xص��=O	�O�%X�-k��N|k=Q��l�m-~��6�H�T[Է�Kf8�8�� �Q7�U�������5 R��W�tl�PNg��'v��X?���῞�~��z�n9�:�yW�(��j�K�!�)Q��w5F�I}Z�[��S�<�#M4�t���[+DoX�aj���^[�Z����Y�������(���]^�1��@_���Ytw`�Hvl���m�4w�����&��F��D�ȑY2+ [����.ʳ`xlk%��yP��c�@�/�x>~����l-j>��,��j޵����99���<�g��4ra��s�٭����n"�Y�*K"p�i��өq�?��\ ������?�%�~�_���������>��'�����~���u���W�O�Z/}��[d����Ҳ�fN�d�;���eVs�ҧ>�����ٯ|��I�.?*����1��9Z���~�����ė��(���AV����S�ڗ,�PD��^�<s�K~Muw�׿�}�;��[ފ������
��R	)S�׬~m���S�Ǚ������_4���ݶ};b�贝�}��=�}7���?�7���Q-,�+x��%}�9�����)|�S_����/�ُ�?Oa�0m��@ �Xgw�܉��i�|�eV��5��v&`$W�Vq��\�t���{��F�`�8~���p��E�/���0v�؄u=�I�����ֳ�<�X��^9r�����|���'�q��""�8ۭX���lj��ݍCx�5� G~=��$X[PJ���<(��|�����j�I0ސ���6�UM��f�Z��百���g'q��,��M$	`	*�n5���`��_[J8��j��<�X�k����;���Su�7x�����Y�@Aa3�R�=���Z� �4Xd�2�v�9R��ס��|[���zmA�G$����[������_ԎK��/�D[���}L'y�>]�,#y�s�}�hi ;J�0�4C�r��Ml��iEr��x�6)����`A���$xl��ӯUy0{�
�Ɉ��UTW&�*h��4M^jڹE�������������S@75��x��]���(����$fT��;&�I"�c�兏&Z�ֆ�G<XA� � s�y���MP͛S� 
�Z�ך�Ңr�B2+��K��	b��b�ਇ���A��y�A-���0��#G���
����SGh��!���7��ۧP�&Z7����r�2!�����q4�9���?����|	���ʥ�s��LєvƲae��R������O��_�
�&���w%f7�$?8��\Y��KԦo���S��3�؊rmv��\��*'���S����a�C�p�����*&'�V�R�����������>��أ���x���133���yd��}=Қ~��og��1������ o�����԰Q]�e�A_W�>�^�0ߦ0���J���7��O�����9\[���4��t_��'0ys�e�B$A�� ��k���,�S�9����t�D'��6��\�h	��yX���2�q�TD���ܗ��?�����/�~���;�E��|��&0?5�F��KW/�w��E<�����ع�v�P�B.KRH�����&珸ї�<��3���Xi�z�0�/%�X�#1�c|HA�9(�<l�A9Gsu��*
+5+7��-kb��/�FE��X��J�\{��I���������
����ORY_��݄[k ���� ���6-T�E�|o�����Eo�qL�MQ�i�*o0�w��hw䝧�Ch��������m�a�z� S�t�{�s�8G�8��S�06�������}�&�1�I-6`.���dMk�im�������9?��>~�b�HE��"��O�V��L�±^�2�U��D�C�����ى���E��h�[�s��>�t�Qn$��Bɫ%r���c�i_"�<��xO��"|���Ҋ�Z�P�M�a��)��=cp�#g�O����"��� ��x���Qk2�DkĕS���8�43Pr�aS�H#�u��/��/>
ץI��N�l7__G�m�A��^ @�Ɍ!�R�,�u��>�h���'O����6f�Wr�a�9�A�T�r&��gN��sf)(?�m;Ob>;�1��E�P(��3Vdx}Flw��k6p]��W�		i݇���E5�Yc��g�s�sz=�tx�/}��x�uO"]n���/`uaÃ�Ԭ��v��H��nŦ}�p��^x��x��gp��U*/[X��xK\;kߵ�)��M�V����p(h[���-�,�o�}�����r"��N#i�&���3Gm���v�7����Mش� .N���_�<�f��FH�:�"�/ڒX�B&���K��n֏��a����7����V�<QZYWm�����@<�f����8����C?�x˻���6Y?��<��Oc���]<�c�}_������/��3O�R�8�%�X$���b��B����[��%:���*��2-T}����R{h@����5�>E����J�Iē~Di�!فU�q2_@��Z˭)(Π+�/`�x	 ~���K���,�&`y�iu�%�Ks_L�g}�X���pS��V���|:K�B�R
P�#р�	p��vڮ_qd�Ep$Jlb�V��v�tK3�l�2�K�%J�O�G�O�ջ��������PN�#�+�Ϋʁ��3|K����ξЕ����)���~���k�0�V*�i:_��<fn�
�V2��HF�q�Vk���x��O�{���x��(z ������`מ]عw+�mB�h?���iE�j��H�E�\f�XZ�@����	(�m�h{�@O^ �ę�� �ˮ���	i����G�+��5?ɢ����2�b\A�p�i��4R�#�4V��ΒYKz�����%Y�i]cP��zɑ������ǟB��D��܃L�n��{Ѹ�`�k�mE�5��ff���w(�2j7n���o�����}�"�R������#��)�b~��̟�2�o|�[�vU�l�JޘL�v���ǡ�1o9VVm�ޔ�S���<*E�]��S'�`��%g �$�(�,}"Ε�q\�~��1�flS��<�k�"G-T�s��	Z֏<� �=|?>����ն�;���A+/i��T�݋u�6��O?�O}�S���ؼe����8Y��u�7dU͙�~��}��  _��رK������ԟ�-����׾�1��5��0@+>��!��C�����5��w���g?�eZ?�d��,�G��,~��ܫ�ҙ��;Y�7!7����q�'��4��<�|;��=��׼�	��O�$~����ŏ��/��?��x�;ކn*����Ō�68�O��~�_�
>��Ocjn��w��=�"
5
}�yLּ����e�'��-ŅL�#�HE;��X��*Qqi���,��BN��T
Cli�@���mW:7�b��>l~�q��؀�-\ZE�'Z>L۲��Թ�W�~��9o�C��*L�Աh$�y�J��� ���@�wm��/�U�ji�;|ɬ������(���WM²?���4��(l�;?���$���g
F��h��ޗW��Ky�}�f�����x�L�����Jo�Ƣ�v�	�"�,	�����P��Q-�qvfWnN`e�B�[�����t޸e6mڊ�۷l�]��൏܏�<� {�!���޵��݃��6a����PGY�d�XN1�.���,��/�X�t"p3~u�ٲGJ�f;��$L�֨���N��_���Ƥ+�Y�B��B�F ����w�Z�{�/YQ���O�pr>�s��̐���((bDA0���ED�%��d&�<gΜ�C����{���g�������s/է�޻v�U�V�Pi��Ѵ�͕ �� S10���Nb�8B����I -&Kٶ����ٷ��(�5�c_Ob�'~������_ g���'Q��aB���p1�%�p�M�,l��O�א۶��i"^��<�g8	���:Zpe�'��^�w߂;n�%�v�x�����Ƌ��T/��ku���*4�!�E�߼����}ι8��p�i_�M����r	S'�����p�p�o��3N;Wz4��<��}X��m\��q�_�=H�FKO��2C�H{O�3��2�N�/�~;֭Y`߁Q_P��T�(�`�ҥ���y8��q�i�BG;�C�ŕ�wwR��%�DϬ[J�$�Ҹ�k'`�������id�߸�Z\�p��?��Wl�aj-*5��K()
�+.
e6��Ԇ�����e�~���1'��7a�ZW[��Jlil��%���~/'�k�1TQ/iV� ����*QR]�ʪ
��i*˱n�ć"��.�)�����O\s�����/�i����>�ãH3��c��� �({��-�Q.���01�Ɓ� <-�8y	�����G �@9���<�V_���c*w�1z����Kc�$��J*G�$~J'��c����xl���w�R�P�V}�^V��ֈG��kte����}���u�{)Wvh�")v@'���x�x�dr�x�\PBO�Q*����c:&�W��bO�$.�e^E���O^�y�>�:i��9�*�?G���@�놎�za��g��s�/���x�l�8�K�u�!r*<Y$�Y$�`�X�|OPC$F-����Vlٲ}��H����'\�ć�J�f���6[a��݇���h����܍ֶ~����pɺ�-��އF�-M=X�؃�-QtGɸ�:· �$�e�>���ϑA�yB>I{��0���蝽WC����3|N�'x��;	�� ��a�W�Q��Y�,ַ7�����ȅr/;Yʋ	��c���C(B��,��"�J8�6�Pcu?�8r��ɞ�i2��|7����c�:�+�Q��M!L����$;�V"<mH��O�X����Α)ec���S���;��x����NC�mի�7Ћ���nh¢��1o�Jl�p5���2�����M�(��}��Ռ��'�t"�kjY[7��������=�Z5���V��j�F,{�-��@mr�X���AѰ�?|/6w�����cśO�5��ޢ��#n�8l>�9/O���7��߰z�V֡(����%��u�r�X��{�	<p�-XEXN9�t\r�ש�L6U�.'�t�V�o�6S�{��'���={�w��ϬZ������.�.�O��1��0lX-���>���غ~��v��{��s�cjQ�=	�ukWਣC�(�>��.�ԩSq�i_BE9b$FGt
ކX�������k/�5�o!�RQ�aӦ��1u�(����A���Kx��1����L�y�ʲ�5�6�=
SfN�P \ￅ\�}�KB#RmX�Q
���|
��>.���s�y�0��ݨ?��$V�X�U��2ҫ>���QJ_V^�h�[7��e��p�=�&Nf���Mk��c��C��Q(���#�"��"��?@\���D�����kW��
��YJ�b���GإȊ�3N�:R\Q���^Z����*��g���p��z9��Y�i7�~k)���W뢔��1/sJǼ���Ԓ?3CD�;aS�t�;�g 2LJ�dN�T�.��v�N�AW����v�O*l���e�E��|I��Kf\��Kb@��"�{�b�Cdb�ۻ�rk?��L�ö>�J`QW+;�X�<�E[:��V�������mX�����r;���V7ǰfg[Z��ږ���$:Sh�M�[�6s"� E�3~j��6��Z����Rj��ZE��[���/!3/��g��f�.��\8�l(�$�f�4T��vx5�4
3���?T�M��~�P��#*"iL5��MD�l��:����/���@��Y�w�E�i�)GQ[I<WLDnƑpLTW�,ͺ;��T�ڶ�\��� -Y͖�E����࢐wU��{�p�q�hDǟ��@����G��1�0O7�r�?�xt��c��-hY��Zs���A���7���l2oj�s( *��m��^�SO<�ΎN�3�_y%�?�̟;-�H�5b��Y�6�֤�e���׋�W�'ҏ�;۱�-B�r��c�ŗ}�����"X���F��q3�B%q��e�ܢ㛺(�Ĵ���̯~g��%2�Q�i��z����3p��o'�j{g/y�~�_Ef�?y��n��3�w$�� <��4� �W)iw���Ȱ�~H�o ��R/�J4�u��y����q'�b牽��v��I'�D��h��a�� ���	D�/a��mظ~#��o�L����*#O-o��F�_�ub���X�j1���ox�g0q�~8��H�,�<���|�3_;˘���э��RZ��RѠ�B��B-#���_}7������/��َ�q�,@��Ν��1�j�Z\�[IY-y�!Zzմ�J�;bCرc3v�v"3�ގ������>����|��ET��y��)|��R�Dr!�u�(���^T�, qa�_���E�-���%s�S
f���ֆ��L��J+x�:w�G�]�C&�|�������j&���$tv}�@��	���(��r�(1#��3��q|�O֒S�W��kKqm�8q�.��1:q���ˣ�����ya��h�XD���Pt�)�ѯ�4	J82<�&�5��f!�s!��`��d �'_v#J�'��7R�Ma�?�����,��}Tƀq6^<�G<�f�,�ŧ��r^$]�0he�M˄��G��(t���mW�K�.�#�(T\*ΕĐ�.@N|'�� ��v�u0#�S!�&�����$̃Ǎ�����hYmlk���m���`�{���2n"��l֐I�qb�":�I �,��hv�q7��\U��H����~2�'�=k6�Q�@u6
��d��W�6 2�t���J4i9��(��߃\9ߏ���j'���I����˗ِX/�<�0\y�U8��)tGb��-�QZ]��{�ZvZMH/Y�!��hĔIp�!���ԡ�����u�Hm7L���O|�¯`�^�#.e9�y�L��3��}i���Cl�z<��S$BM^�(�\����GW�N0�dz|����H{Uer�1u��8���p�!s��!c���ä	�pˌ	�5bf"|e�����ѩs�ۧ�~K.�N
���L�<�$���[1j�@a�!��I>��p(D��D��ٰ�h�n_�!�o߂�m���S�ƌ}��EK��FUe%�8�,xЁTR�O�1��]��@Á���61�%K��?z0�f�L�LgQƾ8a�Za{3l�:��)�Ɖg���I�Ӫ�P�[���4-�^l��پ��t[�I�׆��{W_u5�7���v���]�
�����T2�e�H�k��u--�!m�PZ\b�ΎӇ,�ڻ�ѝ"_�Ұ#�O�K��c�)���s1�]@s�:���k�h��'�#�a���}Y5&,���Bĭ�9h���n.a�x�/�/�ps��v,�ZU��/��M�����.�x�����Nd�s]�(�y����կT��d��*�d%*�����i�ќC��.WJ�1��m	-������
}�Ғ�l�����&��4�4zFJ�����-��uҪ� �e��BH�=S���dޠ�'M��%_!fX���p�Ԫʰݴ6\%E���l�&�4�f�"^UKݴ�����~>6�ƒCdڡ:jE�eȖ��eZ}�)#Ik��	~��f�A�ʼ��^�q�䒠�7�0rS\�'$8�������$ؾt��t6#Nm)��P-y$�U��V`lvS>Z���w�*x��%"��eTh�[	�(oo����� �g0�ڏ�޹�Z����V��0���_ĭ	K7����7�R����Y��@�tG<ytT����c���g��[����ᣆ!�
������Dij|[;�B�w�uh�I�ʶ�!G���yg�Z���0��G�:
�ПJb��d� d%�q�A�q�/�"Ue���.��Y8��^��r��j��Wy��`���dY�1�sXU��;�&��i�p�v�x迟s��b������E?�����͟�qc�1u�L�!n��l�� ���L�����iQv�w����ްO<giؾi�m���������|�\��᳼�_�����>�0t��޿܉{��'��lPL#�U�����+����������/=�������#��B�*9��%aD?~dfL�@6�h�o������%_��7��w��|�˩��_9p:�[
�+8���� )�f�����'K����T����]-�i� 1��� �3���"s�34�b�����X�H.C���-\�Ox�U�	�"'C'�$��ԉ�8�*o6,/�:�'��!�G�{W?�wQn�ቕmx�ݭx�5��;��mdD6JG��0�+��aV���U)�����r���GϢ))�U6��8��������{1��ks�$E'\�b�b��jdQ�5ye)�*_w�ӣ��8ސ�*�N�OR�K��!D�)v�	�� ,��+;Z�p ��"��٘�4�%�ie������ ��7/t,{��n��'�® ��b���(���r��0J"�R������">A��4}fpY�4��3��y��]��a��H�ɦ��miJt��5�$�[Z���܄ޮNt�u#�׏Ρj~]Ɛ����h��Y�h�k�R��p��
�&0�8���������e�yX�r�<���ϐH��r�~���k�Yȅ�ؒm�@���<.��˯An��D��0m��ӝ����4�)���>�PV^i
Hq9;"����K�E���Gk4�X2��� "�f�9���W!��:Kk+ƌ��,L�kī�J{AX�Þd�LD��"QEz�>�V�������^I�-�OJc���F��͜�L�/7�v&m�c����L��A�ق,��;����
�v���:{p�����`��e�����Ͷ0#c`�[����q.����W.����&�r��Ї�:�#XD�vӶu���7�`�{l�
r���D�ʎײ���n�Qp
6��j����GW�cO���>�|�=��ϯê��i����R*���
�U(�E&�JX\�v�>jgۦ������Cf/�1C�$q�q�"<��_�;��v4�4���EEE�F��N�88��c�B�P@sN�4aOe5�����餌4��7y��[�s?yDo_�BE9�Q&���)k�}3wQ��4������PO��]p����+��d_[����<���w�uo�o�&�撣 ��ѷ{h�e�b�l��Q?~�υ������v�w$��dݚ�u�����E�!&�%kG}�K>^ɾ;��S��CI�W�Q�d���I?�:n�7`���O4�v�w��y/��<�Y��7&��>&g&ٴ�%!;�����������Y�7��%�b���S����1/�$"��$�p ��r&��1u��vT=���t�Fգ���Rj��/D��i�X��7�r�LXv	RU	�%4�)x�YDc	D�"���"J�|p{��ې�юx��O���|�vv!�ԅ��N6w`�ﲛ:���	�o��!�Ԅ��f�߶Ӿ��OF���H�q�[MZ,>YI��7j-�V��$����Ѷ�⺊���]�O��僖��iEm\�;� O����#׸ Ч��A�3�/��!�P5�d@Ir�
�t��}���(d#�$4��N6NA���#���b�|�!=��[i�Z��ʐ���j+��C���[L�IE���"��E-�`4��@t��4㗸�7B+�ܲ�1H�־e3cJ�	gil^��7�g��3�2�C�zQ1g�)��N���*_��'0�}NC	�Lt�o�o��"n��	�ⲋ��z��/^�~�5)1C�IQ��K�X�f[����&���N8W\�-�L�I��6�݄k����F�X�cƌ×N;5U��8n
֎��'�Kq	�/��wn������pU=y�E��'?��5��6~w��s:	��^�nj�I���	!�x��݊%�^�]��%�<�B\˝hk��o~�;���_��M��N�sz]��[�,ß������QX�>ҭ�]"�g�H�k?U����5j4��N�h���}{�?�� �5ō��Ҹ[��
,@d�s>����+�0�>'m �����A�eʕ�� <��tbC|�>Ɩd�Z�K����3��Eq��z5S�3o������LG�;o0�{����q�d���x2aGii���ˑ�Q�8?�A8G�*�;�&� �M�[��z̈)�G�jQ�CI��W������F�Wh��V���!Z%�nY9�$���DB	-���%x���(bx9��aÇ�z�p�����	Ђ	���Kk&[Rd����SV^��}�L���������4Y<�d=�l��PK������G��u������֌�7�`O�e�t��K��G$w��KA0�܅i�a[l�#s����/��y�p���D&)F/��9�Չ�$}Z#
60qd߾b�ٜ�,Izw6 O�VZ@�����9��*��3
������.%��?� �E@=���j䘏�w��5���.��#�l��M�X�z"��D��>Z8̃O^ %������c:��o�t����ZVQ�w$~�Y�r)v��D�����������쩡R�2�Ee��b��e������gg��[����/<MAO�eD�+�G��u��uׯ�g0�yo����dI�4'8Տ�>�h�u�Ɣ;h����+��%M��(/i�ɾ�K��腏�W�f�+^��;��Fcs�64c��	��W�9s�ͪ�2�=��	��;64�-߻�
\{�8y
�^��������Ӌ.½�ބ7_yk�,GWWԺ��H,���R��^loـ����'��]7\�o~,�r�%��onŦM;QY=�|�Y|��oڧL�t�ֹ1�+��!�&� �<)?�OA�#�DӶjp j
�D������0|L�N�L����s�Ҳ����uRA&K�#A&MK�3�̩�����L�ZM���C�w�n-^�ֲ����++�E�4�	G��Y?8ߺ�H|�C��[����y�y����-G㊿����E|�����?���~y8N��@��i���;��Z:N>���@�B��>_���,�`M��g	Y�J�㽼uU���3�Yb:�;�jף�>�BF\���^8.ŊR�J����C���5}�������9i�� M5���j��J�c�Edx:�f(�D�P�������|$��� �-	+@<dlZͣ%��?|�%�U�"Ʋ��-%�$4��5_$	?	Ae���Y�����%<��zh��C�0	2LX<~7��!LS����1�ʏ�� |~?z��ig2�T�������Z��#�n5�{7M|�þ�C'+�&�TE�$�Ѣ�=;��������<�t�� 1��B�^������d�P��Q�i�J�u��,lr��g9P65D\��SX�t�}[�/�{�<��- t�Çc4��`(̶��˶��O��ޕa<b�0���Q\Z�����������[�?�_^u%zz:1�J�>��}�Ojm�ǽw�gG����w}�8n���x���ĺ��L�ҽ�������T�¤�.�Ə?�G�p"dv��/x��������l ��J}_:1DVB�I1����+C�>=��t΋����W_��O=�ڽ&X-:���OsRjD���Zu:~�|����G�o�p/�G�Ě���������\�/p.<d�{�L���������:�\2�;a���A8�Sq�?ďw^ذ��8��S��μEo��NDYi��kt`�r�pm����o��8�ة\�i��b�dk�i��z���Oi�s:Af�E�}mH��l���>��#�*)H�T��3��_V��\I�O�
~W�.0�p� dE���.)���`��w���
��GO��/?���L^��o�{ n�l&n��4�x�,���W���3p�9�q�E�������Λ�x9+��B��No�P=ux~d(�X���x1M�<�\���"�#�'���UBH�t*�X���X>
��#��{z>v���`At�h����;i(����MCbCJ ���H�� ;�'�a+>�lm���Ҹ�|e�Y�����
I��!K̏D�L�Y���}�;-ee��H(t�q��v��N���J$�)'�o#�iױ樌a�C�<&���d�.
0/;]��j�qBA�C.S/� ��Dc5�tEAZ]!/�)tݮj�)A��@�O�&
Z�_{.<1�])P6b�}c�8K����V֓��H��X�.�l�^6�&�ɐ���q�9���lX�8w3?�DYVI5����,'3�Lk��c;�]�W]z-�v����c��1c&N8��;�8��q���S��lg
F�emMN=��(���<���#8��sp�ٗ`��6�t/��q�V&�������?H:�Ф�ͯo�O�����Bo� ~t��زe+c>�]A7����OuN�e�Q[�	���??����s��@�7�|+n��O��÷�Gܐ�dn�F�NM!Ҋߴq�}����{�n򔩸��?�Yg����"���3����Re�`�����&O�����_}
��>��r.��2TQ)�>����Ї�p�����{���K��xhA7�mD�5�|:~����W�Ɔ�;p߃w�̓O���ط�S~u�
xr肽���̱N�W2�dB��Q��ה����c��9xc>��:�k��Ux��7�拏a��e��7ļEUTVه��l*_:9E��$y��G�!a:���*ƌ�AńY	2.�_�-�ŗ'���X���P(�u:uuf��o�v0Μ\�I!��:���auTf+x_�ϡ��*�*��2��r*ч����_9g������'/��+q@D��.�2��7$�+��Ě�3O���I95Q��[���9���N�-���d���bt, �Nck���S���dB����i�$�)"PÙ�)lX;��dTC" "4�e��O��Qxfd~'�!�d(X��W�߅��"�Ք!@�'&���v���5um��Ĳ$LZFڡM�i�hF'h_O)����f��4��%!VUWu���@]%<�5@M%����_S��F�S>���A��!\�E	1����։�N<ؽ9K]X�G�GWcC���UUۗ0j�J�����:X#���͎@��! 43��=�a��jX�1j��i��� &	�~$�'#[���ɧ;�7�%��2���cCX@�P��u���U8��_Fum��Ø��ԇɳ@U�p
�,�K��7���;v:�	jN:2:@����o�5~􋟡��x'X�]=x��ר9�\f��O�?�ο�8��߰2��	��j�1��1:n������T�T%��']~�~����k��)�R�۽O����u?���<��x������/�5
�G��3�����W_�[�t3��8�S�����lUaEi	�밁�Z�g;Ae����R��l�����#�p�Q��o\�?��f,^���6���+�ċ�ぇ_$�O�����㏿�W�^�Ek��aG�]�.~~�p�qb԰Z�a۳R��\�]8�uO��09�9>��_�C���-�G�������/�v��"�=Tv�Y�`I%r�b�|%Th�ԥ�.1;Z;qO}� )bR8���>�Zg���^B^ά�|�#��K#Z�F*��W`�#q�i{����sD3EC�Z�[�m�Q4�`�w��?-]h�C�>a!�Ņc�����1����ц��,#/ĝO}�aB�p�[ł�^���	|=��hDF������W,ːuL���76w��w�����2#ȿQ���b�Y ���	��x2�hG?��8J���/���
��f\����4w�K�E�K�Ea+*��(���NȰ�5���@Ac;<�6TPZ���(��C}k,�~mb�w]Z��k�J��u�Gi�}~^}D�����C��A	��u5d���uY|���f� a��hsjp��"�1�'0��g�|�z<��=�D�D�6�F����~�/|�J�O�����V�G�CXm�Kgp�-H��Zl�	�f4�����
�����fh5j�-яL�����	W s�Y�#�Z���]�s�#G��>���y��@� �[N�NM�����ᆭ�ְ������������������G��(`�	_)��+1����SP__M�K��#r�M\�~ڻ��pؽ�M��QZ=G!NpD�C,{���tb쨑9f��)�igK�mC9{���̰��+�6���D:N��d)��p0�,��^-��x��1��wq�?�nK��.�*�6���k�����N3߾�G8���1�����$�h��L�:I,� ҃���v�ceLs�2�ja�<��%O�E#: �-�]JV.'�;�	�>g�BEK�w�n��h���~����4*G�AU�x�j���c��ɨ��(���+�h�"�ܲ�'T�#��P�H<�`�l^�"���=]���&�!��њ��xyI�p��\:�q���ep�p
R�Ju���V{�դp��2'�8�Σ�I^
����9��1�)q򛿥�/\f��[���}�{���;�H���{Bm��7��5��D7㼺f _�����!���7���@���aR�S7�*��d�ZU��qs��=��F�0z�<Y����e;�;:g�+�%��Kl�+�M�7ܰ��/�n�P/k���LTNAd�ib�tJӷs�b����(��i�D���	���J�e�ڹ�|��М�0�4���N�,:�97��)�)���8�N��I�!D)�v�1�&h{R AϦ6de2�[+T�G����0yy9�5HQk���Ol�h{�B�sN2�B3K8Ҭ��2Ĵm��3��ԇFUa��#�7�Èp*]u�t�b�Ys0q��$��F�{6�	�5"����م�;��@jXWdc�tF�7�v��&��k��$q��[�~��/ܓ��.����s�]����#�Df���TV��d�A�����9Yl��'��'+4�S���G`ƴ��6u��k�Zi�j#rc��z��Rj�ΆD��*l��\yN��ӧ`��(�.��Y)��˶&I��E�Ui'h#�V7��U�Z5z�����n{�g�G}>�n�c\'����	�eT�fL��Y���G�����w��t���"�P�_8�t�s�W�+�o~�;8��9�����>`y���8.?�N[(�<��4��9�04'����0�'욃��ɐ�,*�/l.E�ƚߴ{1(�a2b}^ڂT��ϗ���=a� i*&���!�}�EE6#X\e�c��PSS���Z ����Ԉ���]1|4*Ū�fl�m��Dܧ��S�Ng�ѕ�Gg��\A�@aa*P`�)>=X��z�=�j�,`���z�f	�Q�p�(���p�q�1��>���;���c�������.l}/�M�t�S�[�+Ŧ�֡�~4.�bnW;2�؛
cUUw�<ȇ;�_W�������/�;����t��B���d����^6��/h2��3A�8&p��c�؉֠���2%���\�LD�Z`@��jk���!}I%3H0e���w-	"+%U����9mjBG�~2��#�A��a.� �� ����Q���z�HR����w��$���+	Tn{r��5D�'s�Pb6i��h�
�� �zW�G�ęG:�B�eꫧ�O+G(�i��=@��@��}�qtV/��:��Ř� =e�ri�$���"�T���@D�5G����f�uӂ�}|'�jÐ�vF���e$��N���E���Ca�֜�W���HM6�G"�O�K�����;
�a#_�m�%�@0|��>�eZ �������O�@�=3��f���f�!�rK۱�A�G��U:���v���h	�h/��)��Ū3y�o�Įc��m���q=��'ZcB}r�٧C����n���y�ۃ���%׽��>�/��Q��O;�\}9�����ւX�nV�m�Gk6����Ə��v�ј:qZl;a\���q�t�|�)h�~�;&kx5ؔ���tq����O���13��TPP�0���¯=c�.M��m�9N	$�<��l�D�~�sh_�P������'�ZjM�/I^��L������IJ%#�/�	�X���|b0��5���i�Xdj���񱮬�����,YGyЕޚSp�C��Vm.�\h�|���V����P̺�P��5`�7!�(��T"�̘J�ⴽ���g�[E��"���D�����6�ЊT�w�8,<;��@XL>��5�JX3j;�p�M���c�g��[��z����+�y&g���5��@�s��Ȓ��� 'P�rdhe�,�DD� i�I���,����F�q���J�hn2�l��L��S����LӧJ��
���R����SCv�d�,�ὢ�$�P�d�b�ІrɆJ!#�X�$�@������rL�Qȹں�h��@K[�i�D�����9�ڍx[B�硥�����隚��c��u��I�[TW�Se�P9b�Y\�g����+��Mk0[@�owL�a_�ʹ"��f���E��`�xLZ���ŔI���قl�<d�FU�u�7�;�D꺻�=��\�"���U�ئ9~�cYjG��}���!勆!�J��.���82���Ӝ�y�]�,��l���p�\,\�ss��&�Xӱ(:��H_�N^�(�|�L��{'��x'|��V�\�Y�"��*���$~��-�c��R�?m$��6�F����GV�tj3�ѷ�س�	�[�µ�]j��Ư��M-.��L-��}*�����eo����t^Pɰ��O��R�4+�0������/������B�u��+�c��1$�F~e���lR��P0%���b��X^Y�QS&a���(��A��M�-��#�*4$JЕ	1��(�X�UZ����Angs*�٧5��R�ĀmX^�B�1��2���|C�4�w�K��C�qQ��RVQY�)2tT�p��*|i�6����,T���P��J�SX(7��W�bJdƢ�M,>��H_���N�0,��`k���I�m��2U{�4L��Ǝ쑺B�I^�E�MN�	���hʈ��F�Ұ$�ZM˦�ղ���Y�8��%���a�Hh�$�4����.�V"���(LRH�"�2
	"�V��9�¥�a�����$�G�Z���|��x!a�����ٹN�G���5@�ES��߈"�n���I�q�G��Ԉܢm�.jDvU[Z��ъ�;�����m4E6�#��X�|��umpu@�'	���MӚ�iGl��ƌäI�A���[S&!�E��/-WTw��l���	G���+�^v���u��.j�1Z<�&�N!�n�Fx�x��΍�nk��k���?�΀���@%q��Ryf}�l�����s����㿂'��o#���}�n;l�x��P4Jݙ�3�&�4�!ZE���@_����J�����=�KM��0/�3�+g������'�����#�>��V��k��$y�e��fJ���D�
7	'����-'a�-b��]�`Đ�LbB}#�}�f�����6FAG�T��f�'?�,S�T�R��H��HI��e�>�.bf���S��@�ӏ�̢S=�sB���xN<(�Hz�m�q�z�y9/#)C%4�Q�h�G�*�$Ӱ�Z�L�RY]��ѬH�V�U!7�@������EAQ^��2���@fX�#JXJ�e�x
 ��"?��,�1��1}Br#��4�i%D\#� �����'�K{O�����6y6bB=*�b�͆�<��(될H�J�PD�!D��OK��IeM��h!�F�t(�L���>j݊����P]K��S@��Xx$�t[�,�F0S(L��Y"w�I�YKD�J��F� Bmc���2�T��X�hr�K�Y�\�<���$���k):C��(Y&�*�p�>w��u5���K1��T�d2m_B���Ϛ0к�4zoڇ���X?�4�~���Q�����qӮR�g+�Ȓ�i(Ԅ������9�t��;�����$iʐwf��뎷�~� �ӌ�k\����WV UUAK����(?(\J40�s��RI����O���c*1b�p�K|К���w��i�N�$-8}�}�)�-1!c(���<��h(�a'�b^�g&�
x�=�:x~���o���+�[�����·uAfʄ�v0M��u�q$�h2�F����_/:�9vo��D5�
?8�8l� @�ڂ���)���/<��w,�8� L-�cbU�?��46�|�@�੮�d����/���������kq�!SPEkc��u�m'r�8{_\����ݳ���G�<1�/��c��@[֯�@I[���;�c���EVސ,��?�1���V�J<=��(���]�X>���6�
_�+j1�nFL��|%<%��h'��iHi�Mp���#)@G��r�g�&�M�ED�Xv?3J��-q��h"혋̖�v�X���mQ�i+jX�(����u����/r�q�n�,�Cx�Ň���QV9�}�9�EyyF����z�A/Z;z�e�6��j�z�o���k'�lY��� �\u���+����d�7���(c$��]�w�	����遼��Z$��R�� awC/с��C?�vx%�9
�+5O�EIE��ؾ�	�����ۧ��l*�������p��T��]4_;v4�>}��H��7��۪�J=��}i'���T���9Շ����024�f� �'h�i\�IJ|��2L��؄��1��9�
)�U6Eih$��|O��b6~�#�]�Ae@hd=��o��"s��p,����cΘ*�諧b��!�[Prx.<r*��U��eA���X���|����K.¬ه�*l�4�Q�:cF�̽k+p��Sp��Sq�Y����C�d��J����������3~��g�L
��5��V���E(KE硇<(/)Fi074G���t�j��~

iIa6h(�@��P^�M{It>�na#�@tT���q{:	�FC|i\W�]�Y�z���~�{�oy�,'+�w�o���L�h=��W-L����F��k���-HQ��1|,݄�JSy$Yk������s��w�!�:�[C�L�&�CA�'BiI9�ETP3i$���/���z�s�z�m�bgW
�CC�>g��,*2O}�ńP����
��Ѱ����ǆ��m1���,q�ڱ )�66Ǘ����F�`�zF�fL)���ӧ�¿���|<~s����A#ii~>���=�=|��!k���R�^�x2�1�|4_��?v5 �>�e��S�	P'��cAs�̝9�3ʓi4Gh��*��K���b�L�IlMlk��Б�Z��h^�زr�;n����<��KЇ�fM������#G`���|�I8	t7�K��	��՘���D���V���Z����: x�p��M�O h�L.�Eհ�T���kl�¥��$�LB�>��l�
?֩�ȋʚ�ua�k���ꮮ@NK��ʑ]��8�I5(��Biy<�b�N�
�_Dx|�ѱ�H�b\t�(-8����)���9�K+��MҹS�;�<��7�{�pu0�!Z2Zp�p��ps1,[S��QS���%7�uЉ���u��4��F�N	L�����&��t����J'(8����5�i�V��|~?�R:ɰ=�4�,�( �����=]�.���QVTF�J����L⩔B�ε x�¡�����|�	"Ϳx��6a��x�r�p�A1	-PH�ڗ�os��p;^��	=�'��+�����[.��5
e�A#)�D�����_���L�(�-=M�:y���s�6�w�F��8���P'���N�"|���Y3٪j|P��@�ɮa;�қ�u
0�X"ƶ �/P<�Ik�kFP�ųZy�DD�� ��$��l�t�:�P�k�_�MnI�Q@���#$`�)�z>Z�U���%�~�7̐�q����z�x���
f��;	��,�`�!b)�Q�ȡ����0�4����kѲq-�}-�c�����V���.�ܯ�����Zz�-�����U!X_��J�Q8y�a�ˤ��;�|�:4nێH���
6N��j0�,�=N�����g*K�9"��ˑ���p�z��?����@�[�G�[?@���[�n��+�A��Ɯ��S�Z�s��d����s���9��N��m���]��=.j{��,=�3�TC�$SC����
R��ațA�O^t��JnY���pJBa�O2^1[)���Q?�Ư2�x��]��RH��\z�D�&.&O(�RInA �_��Zʄ����X��Y��ۇ�_߀Wo�`,�dև"ƪ�Y6~#��/LS��K"�5����H���L/.\�[�X�����-2#wS5k�e��B/�	1�W��&gð���+L<�W{ȇ��A�0�Fϔ���œ!*@���l#�^R��]�|$�BR�1-�ԋD6���%�$:C4J����b�$��>x���-�D�9@�hR��|�0\�M�鬶���(���di��#kJgZ)�u�����`w�l�#3�˄Z�O�3��e�:��wt��%G�������!I�"���|4=���舞0{��P��FR0��@�w�5��Q���*���>!b\82�r����=���+�F��3A'�#RTk�I���������.�
�W}�k�5��������SSe�J	y����x+[/x
^��Z��\���+�����t�|�l��c���9E81
{<;a�x��~ϰOuz���
���=��W��u�ywv��=���������
�����Sw�9P�s���Oqi1B,�Lx��C���J��!��������1�` �j�������b��P,G�֏�Pb��ehd��G��)���O׏{�����@�%/�9�t'��mp6��;�O��O0M ���>��1lx��<�w<���5�w0��H
��)lo���n�0R�:h ��{��V���.��o��� �nG���2�jb��5�m��?,���/��ѧ]���
4Z�9r����0r���ON2��fl),��)�rnJK��駱̴��! ���7$��^�$��tQ�4,� ���i|��y촑��bE��4�D1%A��4U/�e�<�ϧ�nZN�,*�ډҫ�1
��^4�4bc�vEX�)D"�ŵ����ۣ��1�2�@��Da�"4{;M�'ɹ3�Z5�/q"ͺiݼ�YW����hde){�����XZ��#��h7OҬ.!QU�9k��ċ��{�P��$�Uڄ�㕶��Pq(X�Z�^EX��%T��>ۄ�I�P4��iP���V!�׽�d�amd�"����zg�����OqF���ӝ�`��a׽�l����'ݞ��'��bY��:�lp����Y(-fg#k!l��d?�����㝮�K2^��G��4{�k�{<���s��δ�|?��U�V��r}�J#(>���Ǵ
,�bW�'_H�ɒ�eR	�i��4
e��PT��*��tA�N��I����fQ�X�����/�V�J��S����	���F~D�I�!��R�O��?�S"M	M���?�ts��q����������+�}?��]|��Wp�_����,B�k.��O4������{!�V�6�냟H
�,�)-V}�hW��U��n��p�1&5� ���:�,�` ��P|Td�����Fv���7�E�|��D���$��1E�b�Hs-�����)\��l�;u<6����O��<8vXƗ��0l,'>�DKO'���cF�1���E4��J0&ᤧ��7m��������R��lU-Y\����Yn���P)���k?�C�1?�nG����R������E�֒�wEoQ�SY�':�݀mZ�P����6#��"���_3V�N�T��N��b#[{�=��{u=�EC�ټ�R*��Rz%q���F�)�xN�+����_p".��i� �l��);u�Y�'��dknW:;��q��T+���*��pAJ��!�Q�2u�)�PO�O���;UΡ�+�����'���BG��B��,O���g��x��s�:a��c��K���"!A�>�&O��4���FU2��^}XN'��z"�߰��v*��)�CTDuJ��d�gkz�zz#2���!�N-f���g��O0��<A
�R��5���|R��^J��f�'�r��X��M��o��aG������Ƈ�J��cC�8���°g��_|	Sv���X��q�I{�����7���&!<�� �~�|���dW��T�9���0��~��Fzc"sy�BQH��Hj�I��)�2��gK��fB��5sҡ���S��B�Gb��,�Kz�ϺiչJ���y���y�S!�lCCh�܆�c��:xRd�,z�z��L�b��e��ӏ�����@!�g���c������*���Nl�܀�� �[�~"�ʃұE4�C�'BA�b0��������s��1�9��I{�krO� ��A0X�w��l7�`�o���#���M�)�M�`h J-F�/¦�S�����}S1�KW`B���E�{��k���b�6�XK+8�E�s���	L��*�]^���̏�L;���~��Exv����S� ���39�.�g8�#�g9A�}��R��,�����WN���R��ςR�왏���OjX��EshB��y�N*o�v��<�W�[�����ݧ�]�'�ʲ s�h����SQ|d�Zd@�k
�9%�����<�|¶(@c�R�{����Ӂ�^�(�t�v�w����T�<cv�Qʎ���RZ �+A�U�����J�V�Y~�:!E�p��P�Î��^|��֡���q��3���ē���.:�~�<��C�Ʒ���f��o�.�����҃p�W��o.���~t"����@�}�}S
�S&��F�>iR^2�9��=��z�Rat��)2Ǜ`Q~��Mڂ�qQ-)�$tr��-VfZ�g'3��Za2a+�1���x�4fk9h��s���g_��z�Et%Rx|�<5>ڼ�xҖ*O�<{O��9�Bސ���g��EQQؾC2z���q
�(ap��J��c1�b�^��Y)?������]�����<�\D��Ʋ�/r)�Q����eD����t:�!Z��3%�1��8p���,�,���q沧+0\�µ�v3�O2L��g���:ԣ���<�L�8����0w����ￂwO�k(�iea��#��hO�\�E4�<m�SΦ\ASH�kޫ���Z����6dL<�'ڵ,Iޢ�A��=ݞ��}�ى�'�G�
��v�*OF�׀2]֐�� Gm�O�}�����+?w���,
#&�'�K�@l��F�r�)҄>GrppO��(�6x��u��:�8��EtP�0E�j�l�ґCj`��8Nad��g��+���$�wp;������B�{*��V!�.&�eî�h\�� �U����%8rb {��0����O��p`90�8�҅�h�L�e1�i&���Oc��� Ӱ��hm\�9�N�ov��O��9"W	U9ѨbNX%�*�HJ>��)ϺX�Ux���J�SX!n>�|�6œ�5�#+��u�jK��K:��e�c"�QV�Gkpp �:z�N�B����;h��m�f���>�/��;^]�ֶ>歹��z,as7�t.�@�݃�t�te%�,H0�,
���F&�6H{2�M��c�C�� c_'�9[V\�P8Ĩb9"I���9�!E	��t-l��_z�Nä`�\��(�5U������}�[�6����#0\qf�{�A���g;5ҿ�P>O���E�)�@�e�`�f^���hZڿ�&��0��}TwY���$��,��4����|
jo�����{݉���uQ��rv�w��Nq?�1�b�RAz�a�$�셃�Bu>�Kǩ���
�-�݉Ni�ߖ�pK%��/,��GI~�j�,�9ZT'����A+�B�?	���S\�}쟬L❂&���~J'5D+'�d��8;��X"+�OЋ��0j��dl )O���P%��e��� �P�\����<5��>`�R�O���Ò�+F���+�����q��)|��y���3)��4�A_$����AT����$ߍF�	u�f�.tE�h���7��Ql�J���]	;@���ax-`-�%�I)���g�����A�N~(Z�0Z��<���k��>�!�6P6	м��W�N	p��^�Q"�����?Ioi��l�Ǵ�@�UhZP����ѝIa�Nd� �S���X27��X�LSq��S�S��e1��ؐ-"�Q��|�J��]�xn�f;�\�H^"�$@Ii��X���T_T�R���Aum�Q�v԰:TVV0�HR�I�l��;+�<�(ݩ^:�����&��ɘcI
�l
�8R4ţ�.4�1F`��$Z�GgUeޟ��df���9
̯��
�q�s�9�(�ZC_�5��NnI䔇x��!�r�U#�|��㓺�|���Yi��	:7�.��)W��)��A,�Q�D]8�K���9�-Y7��(>�4��$��j���
���
+�[B��u�m2G���ԳAN��L���e�]����~D�1Z�B��w��Bك��H7N�ݰ}�>���fbs��KI��Y�0��&�g�R
�v8J��kg~NC��ǡn�l���a�僿�E�U��k^\˕�<U�1Qy�����a�;�N����y�ه���d��l_ �$+��g%lᑟ�D� ��F�)|��w<�x|���|������%Zd4�x��������q�o�������ny%�� �ȃ+�B��K�m����/�aX�n��Y|bn���=:Q5��-Ti唟y�2���ܮ�����^IzZb'_sB��T��(�y��K"9�N�S���܇�xԆ�4��q�ʊR��>æUR��	8HwQH��*�	Z^U���= I��c#E(�7� �"�b�jJ�ɨ�#q�I'c�t���lnhA�UK �`�����PUYm��)C,#C��ğ�!��~W''R��Y+B��.��J��&�c���5�W%M�8�Ҳpj)Y�;N��T�|:�6�*�β:ݦXv���aZN���g0�����ՁΎ&�5�@k�64mۈW�a�Ztw��RpJ��#�k�aGs#����W�����4�����b��jGӦhټ���ہ�p�w�}����������a�l�ݎB1��%������_I�3��b�����m���-�s�}�Ex-�� X>��Dm�@ܾ��x���t�"���S8��H�8Ձv-F�����=�Gx��,�ۚ�F���T�����裏bӦMV�w{v����ԟ�;��
��t騾����";�D�὞�}�G'���>��n"BAE��?P�C��ڔF�
v��FFmmBF�6)8��o-\��Tq#4�N]���4�$O�%~gG�:��a
O/�Ј�ri���u]x�������=�����o?؄���m7�Z�ʚ���x��x��kp�-p��;�W6����K+q	�W��)����)ŮN=xOխ�������ḀhՍa&�O3g��x#w�����Ӽ�)W��HL�����L�J�^�,����$�X��7�������a�R�+�^�ӎ<��X(��l*��Y`�8PAnT�U�ģN�1�O�(�3A�aT�y��~����?
����13k2���Z�����A�|5lx-��FM�Y�,T��7��i�ih/�ze�`��!��z���Q`VR�wg|��%3��.�K�;�B��K��$�T�I/��Ħ�7&x�lތMkV!0XF#��v��ʕ����S{�3�
h�������[n�~��_����?��Ǹ�����&������SO#J�l�����,�86�)?��c��q�Eg��K����t��&z)�T�CHN:*'�;��~�EH-l�����������wΙ�{o�V-D��@f�e�ˇs����N<�u����9
e*=6m��ߺ�w|�!�����v��o*B�>�H⣏>����g�T�w�Y���~���{�p��O�\{
��;���	����܈�_�u\|��q͏��c�߇�[7#cV
]��Ҟ����.�w��C��_��~��y:�)D-�n���������
.��[x�ч�h�޹~��5���(=�dP����EE��K(�B���#4��x1�-k7b��0�i+Jr1���ӷ�hW��׆vJ�I /�uQ�,.>����V��x�����W�N���^�ְSK�;yg�m�����!�r��M^4R���#dyH.%�ã/tǑ����cms�Й�a^Y:�2�Q�T�.�Շ��V���%��,�����"Y+SȜr,����2Q��\�ud�x4v�J��5�d ��!��*Y�N^�	�\$w�9N�h
��v�!����顶Aym%FN��S]Aka�{�xY��PQy2Tw*�����8\63'��?{{K+�b	�t���	k�0�n���Y�HM���`�Flں�H��s�v|�h!v4X��hbx���cb���4}����B��A^RB��*� D�Wr�엤��BN,���|-ǖY/Dm�j"�����"���(�x�a�����Ob�L�1�%H]���^�O��K�y�����?1������?ކ<�8^{o!�_�mh�ڶ^��ނ՛�	3�U��J㣥Kqǟ���+<��;����x���ُ���ލ��f�7�:�AT�\N�99
1Q)��.����:~s��X����\�����
֯XbXie77�h�<���s��waٲ�|��5.��aV�Zi�>�"�|/甩�'����Y���o�ӟ���/�WS�ґ��ᆝ�˭�c���6,�<��9)k�'9�w����o�}�x�ʘ�u<�~�q���䝷��m������i�V���G{k;F���������>�,�C�7V{���h���
���[������N�n��1d]��u����H�B�*Υ���Z4\����p��(.�DUM-�+���{��[���SѤN�l�< I~�L�w���/Ps)�.�&T�G9g�U���/l��a�?v7���QT�P�OO����z#
��H.�?�j8�y�}id��M�1m��+��r��,4ٜ6��ꎡ���x��pm@r�B-�f�+_�h������@�LQS�ٷL��^�x�sޥx˷9p��W	�1�y=��P��Ai��3V<
��j�	17�&�T(��&���3�J9�M�$Z;��އ��'�#O>�'��V�Ge�4����g� ���с.�+o����>� ^}�%�Vc߃&�C�cƄa���ƂE������k����_�����'����<";և�͘��Z������� 5�[�z�2� ������$��a�!���&$s�X*�g���7�<���"g�CYG2��� Z�aޒ�0o��2�2�6G�qJSu}�&�_�<�i�l�0}�����U��Ry�hD�bJ��K鼦��x��ǐf�P{XS���i��Au�q��_��{��?�$�{�I<��S��Uנ����#Qmش�ßq������+p�����9�}[;����o«/>�^Z#6d*"wH�~�+k�@#l���+P\Q��}�G��/oƔ�{�%-x�(�7�H-!�cТIa��{&��&ڸ�����_Y�6<�8N��g��}���.���>��F�'?��=�$~r�/����EOG�����&_#����y��;�O�Vz��.�����1�#��Koa���Y̃��M��$0uj�_�r;~������5J����Gww7I�)#CS9A&��{s�_��,g�),j�S���;"�s��N}<�ǖ�A��.Y~?y=�Z0@E74�*�>��H�/�ʢRh_i�y�Y;�@��O�c�ӊЦ?�$���]th�WɅ��;#&�{1j��`H_�?%oцB6z��+I�{{�k]5\GI�+c�"�@/�d�4�E�����$-Zy4HK�!|yɖ3ř0����u8*��]�nW%�Uޛg� ��E����Yoz'��@ɕ��lτ��3YZ9�q[���|
�x͡�`V֎_`�g�2Y�Ȱ�8��GޝÊ��x��7������K�5������)}���ڸo�\�ޞ�g_|�q(���V-[M��B4���2��d�F�[�ϼ�6���Cl#���a�}�-�?�Xo;�oiƢ����[��WޤP{�wz��s��VѦ�4�"ȥ�wǤ.e
k)�S<&��\��1;�r�GHKtS���֞Hu�iP�I@/B��[C�g8���h���X��_�ׅמx�>Z��*�*��8@o2��i$�4��N�W�`��18�S����ч���E��o&���jI�԰X�z.֮^��R|���p叮ġ������_�����4��O�����ټ_N+ I��V�9h5WX	�s�N���k�T#8���q�e���s����9�0��Ѻ%��ϲḻ�d]o۸�GKOX	�/Ų�K���������n@�<��aI�k``�aL�1���e̚1�s�M�����}�+Ku�Y�N�RF
�ӳ4�z�{�`���8��#1�yM�9�~Z�rX�r����@Ҳ̡�����>�tЁA�3c�L��Ex{��ؾ��lJ��ۏeKV`͆��N9԰�>��x����>w��L����eE+�q�h�٧�8|��gyL4:h�^��`JsW��&�����6��:+�Q���䴛S��B�,�\���X�_5�xJ�(�@�ʪ��@V�ڄ���I@zg��(��Re�Rp)ӄ�|��{�S˾"��wx�WF�:2y�)��h��)��L$<��Y�t#|�oJt|~��Ni
�����=��~O/8��}L�$���M�3�R>If��y�R� ���`��%��Pb ��"����~Z"��s�vd=�!���;����=�}�Ѓ�	l۲��S�D�c�f465S{ފm�Mhlo����0�`O�Y�!�gc��Y�T����@���i�j�jlܰ���`XY,���ǰ����	�>�����"���t�Z2�����ŕ�Bso>ڶ�N;���e��D m�/��g8grZ�1�G���'�њ5x����A���Ƈ�(z���AYn���:����A�iV3��8i�&CXIDcR�����w���m�q�a���SNDum�H��U�L��}�L�<��?��/@LL\�0��&���;�NH{-AZ+������j}��"���G�k��ϯ97Kb$f���G���:��٪��ɳhnl��G& ��U�Z�	c�+ G	 D�j�����/\Z���ZۗU
#\T���ؼv=�4�#�#!�tΆT�M/��q%�J$���1e�d��Ĵ�?\T/����62�!2MZ'i���4��g��N-_A����n�a�&�Ǝ�^����IU�1k,�D�TsG}�>�i��A���me���!�u�P��45�����1������l��BI�*�@�̣q7|����v4���)ҭQ^��Y��#iЄ������w|��ov �z��n�=ѷ�V���>�x�*����{ҮV�)�Ԥ�����{�B`l0��t�p����8就dg�HAE��xy6���H��+_��=��4?�IS �*}�O��I`}1_o���|���G+T�!�@��ʹ�}���J�bi�"��{�Z4NmUc�U�Y��Hw�dj�Sp��3�﬉p����]�f����CGs��k�k2�0��&MM�Tv=�x�yx����)r�}'a��1�2u"�����gMe1FIfBpD)�ڿ���EEi�ꆡnx|��:qb*:�)��Z�KMĞ�T��'��9KB�yL�����~��ԕҁ�Ԏ�L�X��:vO��>ˉѫe����#T������Q@$bdf|��x�5 ��_v.24}�71Ѓ�-����K멗����?J���	N�-m����fΜ�q�3/����}�٘	cPRYf��cg�m�C�9+�uU�l7����%:ǅޛ���v���X���𧣦��b����خ�Z����f*!�i2���F������"��RApA�\��3��d��XA�,G�,���OŃ��v4b��5�ţ�/���G4�s�?��:Ǩlix����dBE��&#�'A�(l4ߩ��D{z{L�fG���`��Q]Z;�m�Q��^S���p4�����ܦuS�)��>w��'�⌍�3��iAL*o��S����jٽ�K�L8Mڊ�"�'�����e����7HB��+�W�SK2T��A��E�?��]-*��W������Ͽ�w���TEHh�>�6Ix���o�Ҭ�)D"q���p��J��O'���¾W�~r�����Ž1U[&�� ��ū���!3#m��U��-o���O{!ͳc�yB�����N]�8�ܮg'U�g{�>ײa��\�f.e�.}�NO�b�ӝ��Fw��2�t�Lؾ8d�}p��c���`�0�!����;���p�	�����ч��= ���'N%}�pnQH�H�3����O9g�p8N8�0Tԏ����nmG���-}K���9�pΩ�����'�Î>uÆ�f�8�}e�CHF;��F&#Ҵ���!��e����0��cȦ𡖓#�SB��V�0G���1�wđ��-��ND��|����v$3+
csk7^|�E�[���� �̈��2ۜ�0���4W�y]~4miē�=����;��><|�=�����̣�`ò%��4T'��E��+�5�(.)睆ӄ!YL2�2��ɇ[v���lu�p��K�������XI.<��g���};~����?ބ��Fj��M$�b,���ͅ��`�u�`�%�)���ܱ�9)6;�T�]ǿk�eA�8VϞ�t�J��������qc�Zق>l;	�K�"N��9�*����fg����l#-m׆c}ۅ��%U^F���Aw/�ĳ�2�}g�-*(+/aق���§�
��OGF�!�a�B���a_�C�MŢ�a�Asdd8�Z������DEyn���L"��6*,�)A������~kSF��(��eDe:@뢼�Vm-3 �$h{��n�1�y����Ym*��g8G�²u��f��K�
�	�I�
�J
�{�1Q(�/��:�55�kI�_9p�v�x�k�����/�8���.@$�²����s��jPE��Vc���?'�d]U��� ��[	A�l�g`�L%Tv�aF���tR��[=�e��T	�E�h�m��Z��gm�B����ڝ%ۦ���߸̞2#�����fa��1U[�JZ!�'�������T�8�@�7�����)�L��2H���2��B8��i8���0}�^�k�l��8�B,����ة��$
������}f����aG��,Z]�&�Fe)E�iװ+X�$�0�Gu` ���L��3�aC��h��L6�oc�8�Lu�[��D3��� ��K�^ɷ�sC�;�S�4)�h�n��~�����p�_���{�w����E�b��JU8Lˁ�̎`��ìS T���Z�7^�{\��/�G��7��7ߊ7�~
���;?ph0�t4Ƽ�(&>=T,"/�s(zPS?�p	:Zv"N�$.LLPxh�X*��:6�,������MN�:��ÙT�����������$3���l$��a.9�ZYEfK�[Ma��ք��v,]4߆%�Ѡ����>wH���	Ӭ��N��1����*3��%%����e,�^��h�R�_��ۋ�8������MM[���j�kUX�ʈsL����:�xT����P	+�ۥo�(�d\s	^�b�σ�S��K�L�uhW�r�I�l�P�EH�$�\)�*��ݧ;�9^�+ke��L4����V�����Ḣ�b����N1zr)�^��)aԎʡ�<�}%@iQ�0*�p���s�[�����ӽ=�D�NV�x���\v��E˧��4D�eѼ�e�����+�㑹[����j:�RV~�?��9L U6R��|�l+n��|�����e�iA�t���-�w	:=ӫ^���;SrJ+açBz�Kt�W�}>a�)�eS��֧(AU[}y��,�:c6I�%d�Ym� #MM5A�8�p?5C�+�ظ�FU�����A85�I�e7����'�ˡA��;;�i��\�BSeI �'� TVbC$~Z�C�ijBn�Z8_L�5v�(D!5�~8�K�P˫���e�u4l���\­Uo�6�1�^����{2S�~Xqc���N�Mje��ZO�������XkH�(ʜ�Ći$����g:ÿClI⹹�~^�����
�y$�e��������5�0��IB6���R.�"	���b��q8�S�/���|�]p)N��2L�s4�ť��e��p�ną�3�j2�ݴ&�-STT�)���$�@f�z���r�R,|��{�5,x�ul۸�L�V$iCsF@�$�����������g��?���#���4��9���*5:���P��nĒ%�u�f̟?���&O����F[ԙX"�4�h��ո�{q���ĝw݉g�y
=�]�i��9օభ�����d'�Ҥ7})N%���p�m���[��?�z+{�~Z}������-|
-c���<�h�h�{����BEC�>�l����
���|d�{������gDds��	�/#�}E�1Egŧ�H���b\�?w���>v˾A�Uָ�����Pȏʊb*z%����ͥi*�i*ERB��T�#�8��^�+F8\�7�,�d+�2gs;,W�i��Ȟ�[���pz�wlw��gE�Ւ��jʜ<�^�E��<�V��rCw
�Vu�/�-��o�Ē�hj@kW;I��m=��ҁ���`����x��po%sǴ�Y*S:�ӀQ�ևx�R��3(�'���K�~"K�ra��"Q�_a�"�F�&;X!IT]U�R/0���0 �]�����¯er����
����Տw�_��|}�옑ljhA׎r�$�w�
��lܱ�����}+��gc��DBH�M�K���ln�o���̧ߍ�kס}�T��4��EҠi"'�ر�˖�DoO�\*���|Mr ��2>�9Mm�Yp*l"��g�d�d:�)N�;D�<��9��U��u��+#���"f�:�8����sP��ykO���0
��79��9�t��㕷�a��U���i�G��KQ�K&P_]��z!n�������������Ɵ���^�cO9�>.����U�"\"k��$azZ�����,�i/VU�0��JM�mݴ���f�����\�=������z��L��TU9�6��w�QU^�a�%8�L����	[�X��𞏖����!����e4Q�<�%棃fܘ����1(�y:}x�<�s�=~�_������A�6��U�1�����4�����Z�pސ�!I�
�@0d߃Z�r^z�<��;x�w��Ko��a��͉���l� z�z�j���H}�q*1�U�dl��YF X���
��.�����j�I*h�_(�e��Ib�|i}�:�����Z���6KO#�r�z��OuZ%�KO�C����3}�W����2��iJˍ��5L$�$�n�H���Qe�QU\Gk��(W֒$Bk0YL���[-/Ad`�Mծ�[	{Vk:��O:Ղ[��l-�||6T�]�w�[mkq%���M������Z���g7�O�,ƭO�۞^�۟\��_����9�}!�}�Ʒo�mj������"F"�,� &l�`�B'-���"� �V�'���������ekބ�֯;�n������l�$FԄ1~X5|��;�Mf�8�w_;�v��@_3ZZ��%��!��Ⅻ�}s#��߆��!��I�V ������<
��5Y}b�Y�"-�����H�¦�q���_�⏖ F����Lk`:6���Q
�'���  ��IDATd*N8��d�*�X�
C��*j�(UF��SK�!"ɸu����%/!�H�,T�)���Dr:�=�����K�j��bƼ�:O���Derl�]��<��jjkPU]�Y�fਓOBI�x �j�ġ�>� t��$[���k�t�e��U�����\�E>
qGȉ�*�*QFa$a��҆�.j�7k>�)�z�1�܉T<�a#Ǡ���H�(\
Oq5���-w�8D��GE���Ӫ��Q��Y�3КA*�ʬj�]�Vm�B�~"�E*�)���֡���|/<��a/�p�!?m{t.�A�HeI͜��=�B�x�q��_Ɨ�8u�#�}2k������n� @���'$Y*=	[<"}WQ
��J�ɧ}?��W��ڟ�������Š�rJGׯFw��4��C������vZ����=e�L��a���dh��cm(6�u���2M���L��S�ս���%u�%��s�.�@���O��۩�Qxh�[J_����i�m�M	��di5d��م�=@�-?�RB,o�j/y9*.j�j+�J���%�g��K�$�N��NĪ\I����Fe��!�BE��~<��v��o�;W�OOoÃ�u���q�-x��6`���\ZzNa#&X�\B:z�8� �W�!�B\>� ��d\�m^��@|mY2�Wd����k��jChWQQ��>��)c��#����Ag��ձ��u��X��y�|�N������v���𐑧)L�[;��U��ٱa3�.Y�%K?"�y�=�O�Y��p���������?�����_}O?�֮]�(�M5 	i�B[K;>�p!-Z����W_~s?����n
�,�6�&k$D�QV��Ie~k��e>��, �T7,e%���@Ww?����j�MZT�B��OIӲ���Vf.�G��NsGI
�Ho�{JqW�Yq�Q8���Y-�6�����Po2X5�'�9H��V�X�
��C�R�/�(|��a���6�����X4ۉv�GD#+`Ѽ��ִ�`�6s_T�T[�&����F�q�=���λ����W1�uq3�Zgr��6�^�dr�-����(H&a�;Fc��%���^#J!l��q�k��I�A$3.,]��̼ǟx�(P���K|�o!쁀Gyn������}�x W|�
��5��(�J�|D��X�c�/|��A4�
j޹�F��S'��
PH�0s�d�y�q�_���^���8�G�&���.**�PT\B�z!V�X����Q�پi+�T���F��&qf�f8���x�W�v�
��_�~�Mp>��ì�Lǘ�]�!��&h���<�������}�sp��	�����~%(p��W�v�fca]�>���q�ָ��x�'�����o�H{½V/flJB����=Hay򟄇	'ʞNy�[N�Z#�0�|uN1l�P��u�GD�*�F��r�8���јq�h���2����-�pu�0m�xr�T�{�!8�;���N���G�#;��l���ysV0�|����/�@ϟ�k��Y9�Έ�S7G 9|d�+��Z�b���<I]k�� ge�<���P�t��J�ɍ*��:׍Y�T�`�v��[��X���|���!�}��x��yشq���)F�����������/�+n���a�F��TQk�a$u0����}x�w���ކ[o��{�tw��*TD��Xs��!#�������?������E_o	.Ϊ���܃n�4O�Բ�t<�lb��;:����g#
��&��6��{��)�\��j�	�Au4W �q�%G�K�&'M���^�RCsc���8���P\\��U����,g3feWP[������1�����0�o,�i5)��1�U`���E݈�X�r��A,~�t��@{{�� >p�5l�^{���h�v��J�1���ό	�g�DL�<eeE2XD�VΜ�D �?�V�\���Mx����?���(��wV��c�
P_�}eM=����I�Z]��t$����%̓ɤ�� H��/�.���PZ ��������Z�6n�h���u�&<���x᡻����q�zx�Q����r�o���6���G�Q��X��?q*�\�x�����������#Gb��bҞ�2/G�l���`��v��}x�;��=w؜��g�M�9C����ssR��F����+\��3}�>�	;��G�zn�U�T�}��ґr�Q�x,n'P$T,5''���������[�+�� *����!���6*�K�g�<	;z�P	<k���8��	sR�I�6���*G�<�v{���w�èW����?����ɕG�W����ink�0�.��g�ŏ~v ~s�l��1�������w~p����̙p�z�ޞ��yB�Cf|X��ו./\� �č�P�w���PE��X��t���n�G)��뮿���M�xcYb�l%�V�C9vo*� 5��^
�-+im0-�{��R>��ˇ�2v_jh:S�(�Ց���C�UV���ڻz008����a������B"��e�G�8;�m|~�BD�2�w��A� 	���;�Z�.�G�����}h%��k��th�}"@��OS��8'�J���6��Jp���od	��k"���ټ�.�܄%P��Ec0g�tL�6��&�)�#*�ķ���9m�C�q�G]]���e9v���R�y��HA�m�f�u
5�s�9��|�9j����P� n7c�B��-;�ܴ�����:�J����f����m[�c�j4�2hli��E��|�.��ѓp�5Wᨣ�@P'�(������������o�{�#,[����Jm��Q�1
7�4i�ͅhn���x�V����?E��Qh���>¤���N�������x���K�xA��P���8u�88{K�8�!2��+�b媥��w�jU�M����=~��I�T=Q�\E�N/�OoUf�����fCū����%�QQV�+��=}�aF_a��X�ۢs�-��'�)����J�5�V��Q��8Cpy�a�|�aL�2���7F��d������;�pZ��N��F���÷�U�ȱ(���"� ����_���\� [�����>Z�.���bl��� B�b*$غ�C�Z����H�GZ��)�Y�
���Ź�hʮ��]��6�^Nʥ�4�5�d9T��&T��'���_���'�c�"[���M��胷,�}.���.>��]�)�>��|H�#Y��r?�aj�*�=6�V�|	,2x&a
 n]��:Yf�$d�8�妹I����ty%0/�(罚I#1�o����?nX�ҏז�D<J��g���v��"��&=�d/��PO0dCn
u���Æ
�yki��J��%Ԛ��[{e�H���a�"C�Sk���2ρ(�>��p��̷���y��X�I�.^l����Y��C6g�Ih�D��>����i�r�*L8AF(|t����gu���,�樝c(W��)a�1��=c�)
���k%��+���5Sq��ј0y��1���uw���Nm�+����7�|��d�j�W����J\76�@}U-�p�q8��㌰��4��-���hjm���j?�Ȋ�K��LO;�G��z2;�a�%%6�E[}l��[��;b�'�.L��/�}�wp�)�������m���|u4=�IK����X�U�hmK��pY�۷w`�}��7/�:N?�;Ds(���ߏ
�}���/�*�R�|~
�6��o\���bX]�}T��#�#��Î<�xSy��Id�#���^iImym�*>^Վ��s�ŗ|G�p�RK��W:ej�C�ú2G�K�~��(-�a�l����}�b|���Q��I*]�!�
����)�"}�P=b"N=�b|��`��gي���S��|6j�>�ۤ����W��|�_�Q��{�n$�&�>e�ҊY*���,��D"�Do[)|�S�N���2T�+�J�[;%�J�lm�E��|F�!2��&q���=�h�{��O�2%gO�oc%@���MȖq��q�ɳ�Wuw���[���lC���
�r�����R�=�-�=xv�z��*����GԅQ3��}��v2lףo�c�F���XMs�Xt
6��u1D���2��U����K�'gi��>Y����G6���V|����6�^K롔Ǻ���c�/���=���)Ȝɣ�����A46H���0欙gIDo15s���`
i�e���{(Z��'�3)Z9>})��wI# �>���kŕX�������xZg��ŒZ� NKŨB��`x}d:*�pk�KRߧa~o��ԍg|L+�V�||Б;9[�0�r�&��GO�W�t4Z���S�bG�B��6�;b2ί��Q�{�,o.�ˆ��&�
��/	��9����[�	��1u�4��3��J%iq6��Q�,E��G����+;	s{S�}�u�Y��l;�%�����OWd1m�d�qޙ3i���2	
�n�Z��?��ƆM��:h�8�hL�4a/2� q/���cUS{�)7�j�PVQ�!�}Q�Y�+��DYyx�Mi���0����u�;7m���#Q]Y�,��e�jش��%�0n���j۶��y���0ۜ09����=s-0ܙ���H��m�-з�k�0bX�Zi���\/�V��
�&�g�@ʬw-//)�@]u)�C1���Ӝ%�ۼ���aQ��UVW���4N:5����c�Œ�	waҺ�n����L��Ow��iO���Z7�+�C4���}���޶.��*���~v.���4����՛1w�FDK"�AB#���ƌ��������&�5��j���DG&k�HLU�%���mf�@��Q<��f���{�U<�EGڔ�9��g���2����pɡ#Q�
�����n�������J1�����/�F��y��5M-�텵�`�6s�T\{�^SUas�;�)L��~�>`�_��	��;1Yѿ�V]��F�����!��g������q�Ӷ�b�H�������ET].*��L6���N\�׷���O���Cd)�ہu�Q�3G�30?O �rlo�B/�-�t2.+�����(F��Q P�$���N{K�D��`�9r\Kb�xڑ,�k	���7GP��C�T�k.I'Qkwr�BII5\)&��E�j+�e�����a�d��&x�#d�	����ĩ�!���Ɣ��K�T�c��y���X7=�
6�/�;�գ'��q8w�d>���@�W���V�ut�X�N(��Wk�4�B�%�:SI�>
ksb����E��ND�fX��-<kpF#�_}���֓���r�i��N1g�OP��h)��~��*�ړI��ԶJK���& Y�k�Q|�jO�Ώ�\�J�v�7�I�$�O�*����g��O����)��"��8��OΉ-6���	��[���ީ�*�y��J@0��>�N�
�W�['4<�$ŷ����!�,�h��ǣ�H�R�������d:����a2���ݧ9	t���҅w6��U_�e#�?q������U���c&`��44�c�mx{�J0�5#��&eO�/�N���mBOS�ݝmM��>l1k5����=���m�zԳ�,F�+-y��]�T�5���v�$������&W౫O�i{W#D����M��/c�+��$��|��ᖋ�C��CcwW��6���6����T��:�:}��m�P
uW=��Sm�U��� \A�� �X|F��A���qhS˲%|��<�b��5���L�^�5G��[A���)��ݹ�af#��-1Fpi���/�C��CQ2??���6��dI
vl�(n�eb��=H�H�������{��6��>
'��0L��N<��eғ�	��=X_�=��sՂd��`E� �I���PTT�P8L�*`�+/�>�P�&�%d��bA�$�%�FF'�;+�F���AD��'�Ќ��a�0W�@-������%)3��3�!�L[��u�P���w������O�	Z2F��~�Ki���R�*C��(E]Uj��P_U���R��Bě�R�:ڼ:EΎ)�PYD)q~U���\��=ol�-�s^�iIX*�
qpN}���'\�F7�c�
�L�wrLn
���H�)CF���~��+<8���������6G[6�����/�[p�Z�<�v�[������2�:��u�vU|����0�݋���:>Oψ6<�r��.���	��v2�s��H��2�W�I�r+<k�=e�XP����J�W�o� "I[	륊�E�'C/�OE��jrָ�)��V���Eяm*g}��:o
�u|��/��[�L*hKf>|��+���杽h��I�����>�È�"��^�������Ƿk:�m!�Z܇GWi^�C�n��X�K��ү@�y�ld��)Ͼ�>� cR��
ˇ,z� ����Q�|y_ȏy�'tn�%��$P�[
L�����Hz�1M����j$A�B+5��|Ǒ��9]�X�MRы!/�+<��u�靆���K�$���ּ����I~Z;�t��h�B�Z{^��������Z�B�7��(��J�?x�H
��!b̾��}DY�Gb���س�� �Y�TZ	�"�?�	��Lh!��?�F��&�J�����Sv�DsW��N'�S��T��2{bz16'�Q�p�
5g7��r�"�v��F�:�Yj>�A��YIdg�1�����,�>O��R�ɋН�xe�5-gʟ�m�2����6\���Va���q|4����;=K�:e������>���ݿ��6�� ���7���U�6d'Hg��W+L_��ߣU����>q�L"�J��I�M�Du�>����5[��Α�	J�j^�OЋ�bXa��NtF/�_�\��D�^p>�O���LuQ������1���劆i�՗3S��ãKi�,�i0Rl��$�}(C�)��43����'�NG��	�g'�a���N��?�*c�wz'������Y&Nϳ���r��P1��q��:qȴ>0'ə{^%<�K-ð��a�DԬ>�Pǩ�
E�]Җα������cI�|L��r�F��"YO����q�TZHѯ�š�2���3��`��DM!G�hp0j�0t\��M�L���q�g�>ha/��vw�>�iI0!�L+�pk�� B
D��]
._�^�U��YW坏���!m����)è����+�|_�s& w�Ux�#�f�A��vJ��|��Nl�ɫ���$�@N�ˋ���[�����N�ݠ�����kY��Z=	�#|��,���p�+c;��Kgt��A��E[H�@*S��f�R#/�P%%e|�H�y���!xI�=O�S�i�.*P
�T��|R4�2�"W(�n?������6(~e�d��Z������֑�F<�p�Q�%�0���֣�kz|]���h&� eDh��F���	���̋�P5J���j9�'������TS�������_w��X2'?�N�U�Ɇ��w���1!���K���E��Ӓٓ���3�H \A�؎�< �u,!�Nr�(��:W� �g�H H�h8Niw	�� �FϊX.ָ�	t��*h�R<gә��?��A�@�-��=�Fa�b�=���Ϥ��me����i需�t�S8p����"j`y"��ԭy'�:�ƑY#����Bj���V��a�6�/fd�\ ls�8P�#5��
e~�1����/oN]Ai�iy�ͭ��;r�s��������N�XʝW¦'�κ���3�<��4j�X	� Ly�'7۔��#�dB�G�솯�l~��!���ݿ�c;Yb3��H�h�t�4T"�P�h�&y���*��U����|�	��J��F�Ӽk"���0we��N���a�y�(O������ȍ����ܵ"��Ѿ)��Wư�T���j��,���ž'̂����(���5�4��|�I?����ZC�0&�2�7����G�
f�C�0�N���.^Rp{VF�X���x��C�r*�?�qψ0�%|y~e�"�ſS� ��<��j:�T�r�:�Ŀ���L#`|�Y�̴ ��m�2r����#���\�N1�N�W��c�z.�U�0V��g�ͫl���V	�|��*�a���W=	�.-�7c�E-'�D,1DӜ>�I}'\�*2C��T��|���Ը���
�0k�Dd���om| ߐ��{:v.�O�*ӽ�lW��^pE���L߀�`7�TC_���s^M(���"146lÆ�k�c�6h��Yw{���_�E��uuw!E�Oo
.�fimo���+�q�JD�VGC��5FQ{� IG��MX�t)6n܀H��`b��?QL�R=>Z��罇�;6�*:��ql�9ۭ�x��}�4nX�z��߬��l�i$<m'�o��W�/>x6,�O��?_�S]�p�����Ѵs'�q���7u�|�]u���-�tl ��j��F���Jc(A���i§��J+��E B�K����!ՐV�PJ���Es�A���}��]N��9�؟�;�D<WL�w	�u{�Q{��)i�ư�S��܃�J�:�5����8��^�.>c6�C�a,5�ɠ=2�,��Ŕ/L�������)�Z��-�������`��,����	^0�jb�
�X��"��$���3^O�S%�-���믿ayc7^_���r^"C��&��Isg�w#�Eie��=���F_��Y��6,��e�p��tV/�g<	�]�^Q�F�R5�N5tU��1G	K=Y~����Y��ZΜʤH<N�I2�t�k���&���6��bL]5F�fV����9	��3af�<��N��	�P9��TO���ܺ��0��$z����s�V~c����'�v�
�X� �e(.*e^*�fW�F���/ᑇƒ��E���$*/�Ԑ�:Ɵy�$������/����o����#I&\UU�P�:���[�6mބ�?�[m�>��he*_���㯷ߎ_x�ϝ���+P=li�ƱL�V�b�r���K/���b��e;v,�&0�&n�غu~���2��޻�`Uyy1�f�~�����x���p�m�᝷�ƆeK�����ɓ�-�p�G��e?t�]x����{�`��M��|����#�V�\�Gzؾz9i򤏷����ˉ=�e��x/���Ջ'��wԍ�Ge�h#�>�RTB��Q���� zgW�;����Q��a��j*��
��B�P6AZN;���1g��)+���y\a��W'ܞaL#��+M(�����9ў^��*b�kt�e����XW�ʀ��|�5�s���բ"�䳣#�?>���T��yp퍧�CFهed��с��]��+z��ه�,;�2x���������j�]�j�jr9"�
kV�0��a&�m�E=T����K8�gT/Z�>m������V+ᣱ���4�<	x������_R�T���cYZ�������CĸdT��	�$L�Ǒ���WE�s�*�+%i J�LV1/���	+SK$L�P�`����>��<j/5�4p���LS[�_�_B�/��l�ѣk͌_�O���=�@Q=�S�q�fc�^3Y�p�3�Ep���YNZ��������������D�|�r5B�(��L@0��ʉ$w�h�?�/?�	Ѝ)h������(�}�y���[0�ݹرf3�/]nG����9a�-ʈ�Sx���q'��+����.�Y��V��o�7E%j���R�ޛ��p�w��{�AmEf�5�"a�V����������^�\�==Q,�����|�}n@�hkO?��*<��cشi3z�����o@�P?���l����\�?�~s�o�sg���͛�3�&L7�G�d~.�����_߄�,w�ȱh�يՋ>���?��}l��L��}���W_G�r8*FM���[��т�f��p2#aZ.�L�zیG��O<���()
���BiY������s����6!K�s������W��CE��3n��t��1��QUu"�;���;�Z���*�p�׹Ũ�cr�hݕ���GާM�t�9b;�I�[�`�?������W��k���/[=��M������
�Y��=�AK,�q�a��,E�uY ���(�������-���-T���E��e�`L�҈��؁{�Z�G��W'�"�3�dj�rĿT��+8��:�"+L/$txo����R�P��A�X]$�x1&�<�����J�P�h;�ig��u��K�i֕��0*-)'l>$�����܋��ňdi1�&�yK�R�tZyaBD	�.aSE�Sͬt���-��T&�ҭ�>������ϋc"ۍ%���4�(�7��
�نޘ	"�-���YXNbd���m��&�W�@���x������$^{�<��舧q���|�4<�܋��|����Q0z�E����/�Ͼ��X���� �d�D�.G��}���������O=\~�)H�#s�g�ܰ������[o��EK�`���q�e��O?-}���a��e�f\�m޴w�Ik���y�l�a�#��R��l��d:)�����/�6���cO�y��P���l�Z<���D��N����A���x��j�
ß���=��_{�V4~������š��7�x���~[m),��Y86�Y�#?W]�S�z��єv� ��� ���c��x��WQQ7�������ǟ~B%�h>O-C�צ�6<��3x�g��J�#:�2�Ru��;���U4�z������hIJ��1��+O��S�hZ����l��(���ϻʰ��nW$�����X�½���;�N�|�B��-�b�9_.� ��0��T"MU����k����V�2�����H҉^���9}�-���g2įde胁Y�Q	&��$O��(�"^'XM��6�'��=V��L<#_7��N�MV��!L�j��F�6-2�?@u�B@Æƒ�u�~sK���ϯ���T��"�J K���cK'~��
��%�m��DV��fOg�"��ޏ��Z����w;�հb����� ����U=���+��u�~�6�7{$Kȝ6W��ߜ��΢'��`%ˬ��Bfޅy?���(�2"��o(Xd��h�Wdݨ�$h�@��!*�lֆ�tn��5�H��ڿ��,�J4�y�|�>/A�s���<�>�T  sD����������n4�J�+o��*7��!ل����Bn�m��q�Fl�rԀ4�%bW!�D`��>�鴇�;v���Nǵ��?��z��oc���ݥp�CA��99�N����o��:�o߁A6XK���
О�^T��⢋/��~z.��8��c1H��-[�M��Rd�Y�r�����~��
��կaIX�n#֬[����c��$ܻ���}:;������;yvp�ج��P�Qإ�_���>j,[;hkռ_i��:������]���pλ�|L�>�V*��Ƶ��{`0���(	qʉGa�����)1�bނ���6B����`}}=�;�\:�`�9� 7�75aۦ�*؆�֭]E��ch9x྘:q,N��	8���i!M'?p�����-X0!������M������N?�0y:m���>��'UY�aT�T%)�X����N�3a�g�Y�UY�Hve�|��l���+8�+7�s�� ��U��^��J!��HX<'��)�`�4�yP
�{������ecl��t���>ݑZ��(�>�T��| h���AE��;�7��0�&I�?(���0�B��hԔ1��������/��S�+o���1*G�(y����$9�TZeړ
��rkBT�H2�\7�սx��&���r��奸��������yx�5h{���%I�����s�񷗖��O/�#onG�f*���0�R��m��	�^�r�a����VG�0����mZ��]霴�8^�ȍ��FDrRl'a֕BOo?�6lGR��I�4թ�.;�ۘ6˵�.i�g�����<-��*8m.՞����:�[>�a�;i��
Wa�����$�r�"x���W�
T��J4���Z=GLKp��rʱD�ϧ��w:n\sGZ��̳�$z���j�XZIf7*S�|ö������T�?�\}�58����a�0a�X��w_;qw冭�J�P`�x$����>�7��W� >�><i�X|���ŗ]��3���������ׅ~zկ��g�{.~���ēO�O!��T�y��$�����A���'N���r�ֲTqd"�~�+
��$�r��b�����c�0a08��g��u?�?��j�_jز��1�B::��� &��DZ�a��۷���U���0iL=[К,F��?Ⱥ�c�ڰauE1�k*탂�6��c����~�]OW�}ba������a��Iv��� �V5t���GOk��VV[��9���;�~�֜�LFߎ�F�ҢQ����`v�4�V�����؉h��@�`a;������-����3�:�(n��SC�:���y'����exw�@��ذj)7����������G+iW��ݶ�{/����Kh!��� ��CR B��{�Ƹ�ޛlIV�Zm��{�3���/!���&��{�N9s��)3sg֣�����`V^*���V-��e�Q[�]�ހQ_0�=��r�gX�����m;7+�Dqt�K4��
�?#���T���=�T���Ů�RBᒂ��Bv��"}��o�����p�.�>�V��(ߋ'�/��~�Ϸ��� ��M,�R�������N<D�ۣO4(|R�12�i��̿��������'~4c���8��"e}ެ���m�����R<��ex��-����0�X���6��[�ċk��kQ]�IXOiCB�|0�R�2>����C?]�N���٣��������xOë�S���/ķQ���TB�>�euU5�UU��#���9��K�߫�l%��2]�<zG����G�j��!f�@{�z�>ߢ��4�EM3�p�ڦm7�H��p�H��4��~+ԏZ#�fgLԥW����(b�r�S=�S�I"�	<jAڙA�4l����Lo�����+���#<�tfN�������L�QsSʹ4���6�Yk�$�n֡r�|��G(�S�j��H�#ӊ�퀲ޘ1s�P��HME�VA'��̫d�0�����f��f��#�D������tv��O��)�)%S>��p�7�ODn^�}� ��o�����F������~�Z��4f$�dʄ�wIƌ���l,��#��_��m7Ed¤�Lo䈼�LL7Ά^{�]����Go��<����G��`G%�h�+�HSll
dR@񾽞�t�j��v��v2��Ț5l.�w��ܷ^����5Q1"����;���w0d�cR����Ds��!� k������܀/>zM{+)\D�j�퓸pާx�����[n�Go��:;oI�P@ѷ[��k���܈_�y����l�Z�qZ��x����n����=V��%���Ԉ�A���c��ӛp�ͷ��߃��aʺfFj��ꫯ�f����[��C�|�&��t�56��"�[o�n��gx�Ϡ�v�����U?9C����/�qvؖ�n��T4t��.~Z>ZZm���|.F���t�ئ�������a>ڍ?H�/������'������9�[�F�-�<�2
�T
�T)���%�d��#S���0":X������)5ʴAƓ���>^��P����9٨�"�3�|GFlJ10V;���]G����������#�B��iT��[�a�Ѣ��yz�wa��k��UuJ@'~��n���p��U
m�O6��bggD&T��nԳ�v0<L��&RlL�M�	��%
Q�s�qV�^�CS����P*Fք���
]mH�ND#gK�{�9��&�t\�e��"�!Q{���L�$��=�|��{�D��`k
I�^��,����B�$-��g�CW�6�t�ְ�ʑ �WNy�o[���Zέ��%�#� '{��\Gg/]�5k���#��C#�V���a�&;�!Q�&�vlߎ�ֱZ)>� ����_��vjl���b۷mŌ�0a�x�1�0���q,w�99:��i�ح�a��������YL�1?)#�FA�N2�\
Y�M��X<1>��s�'�C�v�6mv [)-2u�5�w��w>Ď�]H���w�>���7U?���ϛ�t��N���D<Hk��՝oD������L��7������?�46�^b�}0��,?�덉���*�N
򰶌���Q�h�Q��y��7������w�����7�/כ�
Z���Ï���_ģO>���{?>�u�S�5:�>�;w�
�ǟ}O=�<}�iT�qC���d`�ʥx�����K��'���>�9<m��l���_�M��-����x��W�������p"�Q[S��s��>��|���z�m��m�*��ڨ�[�Ͽ���>��w>]��~֭�E?̂����}[c ������))'���l�7���Yuƕ�㳿h�Y}���%�k�����G�YFH?!�s�x���Ψ�0kHu��ū�W��[
0�`��Ԅ6�&-��F�h(Ύv��nڄ3��gf�C�z����������=�_w8����t$���P\����}]}8�0X�@wk�F
S
b�i���(H�q`�+�>���eW��1M�b������3C�j_9�j�Y84F�H�s�VM�e���Ű�/ ��=��yd�1�J���	�Jg��%���� $�˄���$Pd,J���m�*�TiT��˛�g�k�D[ ��Y���Rc�)��Y��z� �;fBX�xo�a%�����F�1o�`����M���Gg�<�j�m����(����:{�<5����hk��t��=�k1u�DL���OC�6o�����i��o��ه�2Q�%��œ�'V}$���T>���ż�<�`�x��dڽ	 ۂ>YǶ�V|����~YY���oc��	�T"Jg ��)�d�i�6$�B{\e�n��WЙ�����<זl/Z��7��4j�4��\6&M��ˮ�>f�:]�ǜ�YG�B���vnmk�����Ob����yr3����hm�kG�t�^t�F�`但	ԡ��.?Kc���1����
��߱�p�������FO����j1�2�:: 酨f�E�9��S�hkm���E���8cf��9����^�v3�n����8.X����k�_�ܵm'>��S�Sk�$CZ�j#�}�IZ����Q@o߲+֮���
�y�޲5uM�x�ؑp�mT�=�@(�����&)·��Ϫi�@��q�x�d�:�Ll'˯��
uuՆ�ڳ���Þ];��"����Д�ql�e�t�b�P@I(h��8U^�}�D�~��q�hW�Td��ڋ�Z�T>��t~�b!�D��^�;:��Oo 	.#����H�������CTO�	s�r�?�{��a7�Qy�ţe�)���	OZ��X;�kOMm��t�K'�@������A'Õ����8�>�6�:7���)}��qӱ#q�i�p嵇b�%�2v�CZ3%��w��U~w�J��r�1����pHo��z�{E�e��o�[3$޻S	�|�+su��&PD0�" m�����d ��|�o{��@�=�%=��"o+�++i^V��U)8�sA�Pӷ"�6u���M�z->���$p���G�&�I� w�R�'0T)�����p�gYu6Y�wI,��I`�=�(�>�����i�ـ?�D�F���4j���1�~�St@̠����[�|)JJKq�w��j�*���s>����̣e�e�}hok%L�d��h��pN0���6|���x�g����_`���#:ˠE�oي�x��Wl�1��f�:Z1�PC��:;�g�g�����I��ꕫl#�ou$���j����*
���b,��jsԾ���<b�-���g�G�]��}1���}M���>NM�	-0�3q�UW�� ^q)Ǝ��%�Va��ĲӪ�i�����jՁ"�(�[����*�7KH�/i��^}�0}�a3r.ðI��)B�{�V0�����CEZ=Ґ���8QF��!���o��E�a�ʅ�2��{O9֮Y��v	G��j���X�t���i�Rx�\N��>:Kȏ1T`���%�'R��v�-�7%�}4��ޮ�Rf�y��TSVyݱv#>y��^�K���Ǵ��Q�)~��ld���kX0�c��������w�8L��6}�*vmAGS������Jd�&���s�:2oV"#ށ���Ho]&�ٖ~tP�
�ڈ�1*=���-�7����څς_B���D�Ty9&��z��g�q��,�>By1]
��D[��1��{��4���8!� ai�3i|�A%��܃0{L/���j?-�xmu�P@�}@If���pƁ��U30�!�e &u���P�td6XT�G��[|�g��z�钸5'�_��m'���V8s�L�N���� @�J�̌�4�mNB���3o�I�U֧/�B��G�F�M�9��H�-��N���T���I~��mb*��d��i�./i�f�(_vJ۶��U�v��IW�:����LT�*�<U�!3���^Π�#���l���E>9FS[�K+М�� Re�A�Ӽ(��Cz�*�q��9��:$*�e��*���a���S<��k�*.�W~�gϖ�N�SPY݈�>��5Ԍw�Ľ�ݏ��x�4GUE�,�Kf�4r�!�Ɗ����/�j�6y�D}�7��IV}<+G�5L�_��>�W|�`)f��8��Pڷ�C�*�:[W�-�����&]�N�+_hy�"ZXbdG5��Ǆ�q'b�YX����C����v���ƐW��!��`�	�+.Ć�[Q��A:��aoX�F��Ɓ�'�O�>5j$F�M�����hդ"�m��Vv��6�9��SS׈�/ː��P����#���TzD�J����T�+���vd��Z�5HL�6i����NZ�C�FlCG�*|��E��h�����x�I���'1��g�E�����I����ES�O��n�����������y�����+��>�jKb��-��R>���Vp��K׺��6O.S��i���/��_�p~s��x慗QUS�l��0�so�x����[q۝w���?BKs�*X�z~q��p��?�̈́��?�5�7���6/�m��vt}O5�0tYQz�#ȊU&FR|�b��$G'k�G�,Z��9)6"�m��18S�5�-���	�x�%�w.\��_4%�((=�>�z��v���V�����ej�7��:�
���%S(�Q#
�+��6¹n�<�����x��(o �v�FA�����"\}�a�r�Ht��v����W�d	j჎7P#)LW�(�n����uխ�m_��Q�\O?�/�Ba3��8�Υ�!ɲr����³<Y>b8&O����<�f��F%m�dM��y{&����wD�<�\Nm&o��H )V�T�-d��f�K��R��i����hR�9�qՔsL"IXGi��氃j�%�`������Y0�"x%[�Η@�ƈ-���)�ӨN]f�X&t���8!�_�t	~��?���^pο�Bd�h��EKO�@�~C1c���v����;-�����^n���*\�ع���*�S+=�`�������vqЋ�(�ݻv�}��.��^z%&N���X!��UKwvaJW?�R�w�Q;!H����#ןA����Fna>����:D���j>��.����#�Z��W�{��^���mV�alX��ۻ�pU�x�P𦙝&EA2~�?���BG{v��F�(���Bd�9�8t�ьv���ɶ�w�._FˈB���UV�z���J�-�p���'����.�1R;�t￲3��.#��-^ͺ�^�W��n���b���G�ȣ�gVa�����+q���}�8���x����Koa��]8l��f!^y��8t�t*�֖�PLLS4n0��#dĲ|I�M�DK�*��[�����h���k��;��\��WbނeX�t�I���:jjj�b��ux���ԋ��׿�>��S*,�6���V�z����t��,�������%���%)ttT��$e)iT&��(�!�H�����$�<�þ�e_w�{8^�Jb-�R�3����n�xji���1a���\%�TO]��
�@��L�H���6ߣy���NÈ~E(
xm�u{�p��K��㝇��;���ֱ`Q٬�'��|/-�I}q鷧`ƹci�77D��]b�K��WL��
���а`Um��\�����ʑ��a�a�U����-%�j�L�s����6ư�t`f���:�S�I��~f:�M�j�|��"���)%�?�*;gu(�l]eL3P���;[vͫ�ZW��KÖy��:vXq���H[;9|'l;mĲ�s7.wW��kvV����*UѽN���FM�KFа��"V�,OKCe[-�]m.Z��	zGp_ꔎ�VUV��ǟĪUk���g˞KK�Z���WV�߹�R�t�m��[�k����W����FM���%�7�4��w��o�Mܤc��a�A:5�tZ���'���>@�pvβ�e��DI�b�r��3�N��,;/�Z�>3ʶ�Y��}4VU"d+���u�rL�p �~?�H{����_��~�;,_�)j���k�f�غ�,�z�2��/(F�aP^݂�>|�M��pټn="�=���ᥥ�����?�6�[��7aoe9��
1b�XBOˇΠ�#���˖.��/>��+�z�b��";z�mţ��9
r�0�98ͧ��L4~-g0�k�n>�Π��J基yc�aK9��؃��F���M�LĔCg`���@kl��*�m%|>|�TL?��K�ZY�nq��o��5�k�pDK���.mϟ�M�o���6�����:xԻo��y��"��$���^LG4ݍ6>o �KV�e���|�,��c�Q\,��=BGS#m:����oA&�N~n�	�s��k�'N��]Ϥ��G<�4)�b��9�)�ʹ�s�N%��%|s�U��3Ho�YT�}ٔq��1�vQ�'?5���Uc� �{K�$s[�Z���ز�ѭ�\��fG��b{6�58
2�cG���E��,ZZ̳��}�JyH4�{`��K�W���g{��aw�T��޸�.,�hw�I4�+AN�cל���Y߼"�h���7�bW���P����"g�N���ʾ!#>��*5	(��iôpi�L�ci�1v$�b\�(,r
OVRs<�0*�c�OsE�&���P�'�4w�z黆h8LSS�+��%�\��x��|}h��I8�W'
1j��Q���F����Đ�S������#�Rd��чx����C�B!l[�s?� ��/��Y1��,?&M�C��㎛���9���e�ܻo4c�	e��ٰa>|�=TR�i��+���ǻ/=�M�!�tt
��*0�9�U^nm�n�B���������\ZBMl�su!yi���9��}z��$�A��Ɋ�M������7�_v�����7��w��1���?�JK
������`�m��7��s/��w܎��V\z�O��<di��3�;�-A�����.�M�\���7���/Ĩqc	U
rY?zz���o�K�����~����}ֹ�[֏`��L�rfy��܍���K������_��I0u�Tks9�Vm$�a[.u�c��q���	��U��> '1�	o}7#�wN/y���)��p&�z��18�>��)�&���H׆�]���	���1O��fx)�����9y�2d�]_���Űa#P�KS�te+�*��,�-������ J��8��	+/���s�w�����tVy�؝~j�������Z��A~a
�rQP�g4,�ҥi��CC�w;�y
.	M�K�P|���;H�U0ɣ��虯t�	2���j��R�y(Q����?i٣�^J�Ce�+!=��,��4�)�-Ua
"<!�:
�X�V{�~�L+��8//ۂ���+�5�]�3�p�B̘2(`fM����,� B��e휊1�`!}	0�	�p��| ���T_��O�'\鵅'�"Z��O���[o_]шV����@��y49��Ai#7քx�^���&�D�hmo��p�������
6��,��*��*��ݽ�c<fSH"�Y=	�<l"܆�,_���)�|��¬��#�q��R�};5�@B�n
�ӭ��$ԩ1�.6�2�d�ۊ��2�,�E��Pۀ�x+�M�iA-�#FNĠ��o	�ut��/u,������g�[��ϩ�i��-X��\l[�'���bC�V�hY��2���C"��O;��������s��@+O�u���Ú5�0�Ӭ��J�eeb�x��m������[��c��5��0v�v�������_�	��8��30|�H�F�^K�3��(�a����;�nތ`S�^�C{�7���&�<�𲑚��O�~F˯�V�.��TS`�g��fg��S��M%3,Bsk'��Y����#���9�b|��s�W�/L)�@"=#u�س����(�}��8��Ӑ���څͣ�n{���frm0ß����瞃�G���d|ѧ�d�xR2p�b��1f�����W�h�,���J��O=��:�c���}[ְ��A{CF���f˗���Ͼ���M6�j�!����"N�Q�mK:Ձb�T/�M����)3p��G⤓N�R3�u��jԂI_y��(��Ç���3	��fL���3�!�L�䃦ࠃ�`��:m&�31�י3ǴC�����0u�a�:]�PL�1��n���㠃��
��I�#f���>�P�)��ݬM��#ވ��PW<�������G��c���x���{�*A>-cm��҆���n��݈XcriRi�����ʻr�{w+Z�jLeIW؉��ܠ�"�&Y[�}����;�ϥ�6��������*�Y��Y� E�vч)}T ���S�b܀l�dV�l�ǯnE��������k�s zg��#.��`3�~q��[0��mț�:ux�XW߂����*P(��acyrH�Π�}�n���K��oF��g�V�E]rV����೥���)-+G��#�u?9�{b��5�;�,:ǋ._�Բ&��<�� M��Yhm��ν{�t_�j/"97wC� & �19`�.)4l���N'��:~a� �O�H�!�x�����J76���\����5~��?���{-�v�mnEcC#餋+��R�E�N��(�f� Q6�v�ѐ[
���`ơ���yg�l�P8��
�a
q��㿅Y�<i^j��(�����5�?v�������7+���VY��[6�O)N<�$�j��jX�J ��ښzTW��С���Om�D
ǰ~�6,�b>��v�����08p"9� �ˋ�=�X�d��*�R���ے�d�Hᓗ�B�^�b/۶����#GF~A.�Fܱ.ڶ=BKy��:|:�47�"��n ����LBaq����W���N������P(�٤�Q��Fq��|�l^B��غc7V,[G"�Ġ�1j�P��T�־����G5�Mغy��0pPo�Ї�-T���&��+�&��N�IJK�QZ\@a'K��y����ii넗)�V�S���p��l��܅�N?K�l&ݫ�h������{�	�˖c�e<���A[[=��V�\��`5��Y�>[6h(�Sq8�ȩ8���P�o�����N
�A�o	���F�J����]̿��WT��n֯��<�S0<	4$JC4��W��1�Z-��	��@\L毓E����8/N���+8��S=Ղ�&�Չ�kV��[NAWK3�d���`��19q<ڃa��U�>Q���6�y+Ѿ�)%�Sr�V:��J0>g�_	-�Du�vt`)���`gK�j5j:�ѭ�U;�C~'z2�V˺��TR�!`⤋<�KR ʖ�J��o%q��"&�p�U���G�@N o�i�e�u�w3�8�?v>u�g(�w��o�埮F��{��Ƶ'�AE���х>ف���	����*@F�l[b���F�ĭ�m�tB�F~l��i�<6ަ�>�vO��~qL ����A>c��aֳ�/�������㧗P�4�l�l�Ӧ�8"��3ۨ�Yd�!��&j�`���M���������7��r	��d	���`�t�6�ԉGBC_�kE�	(��%`4F+m[N��)��_��ؼW��fK�45��v�FSD&�Y�{;S�$�q4�!��%�G^��E ����'!J�q�V�W��;�u��ণN�G�@A=��Y�ܿҌM8�[Z��r�pQb6�L� ;dNBcW8k�D����[�ޅt_��xm������f�C����v���tF"&䕷	L˿���`}��$��J�I� �����Fl�))��&��h��*u� ��<�khV����u�)|�m��O��h��Ŧ��Q���
��4Ҟ0%�NlJP	t��9i�Ot��3<	 �{����)9�f�^����R|?X�,,�E��N�1o]v�ލ+/<��_n�U=�m�w.�^u���;�}��r=�<�H�p��-+�б�6�D�3�Eƍ���G�p�&&�LY�����4*������4����ei�����@R:�W{)�hݲ<����|��N�"J-,�ñNl޴��B4W�ƀ�T\��DZwF��&Z_(�I�SY���|���F��gK��CZ�@2�b�/O��A�-�`Yĳm�M�DV����	�1�RM��+���؅ui���]�9�o��&�L�*�;i#}�����ߜ�BZ7�:�������ۛH��8�ؑ�㙣��c�!^���x��S9/:5����|�PD�Q�w�K�=�)�L.����C/�#ŕ�,�$�)jE���	���b�$|hAh�xU�X��YSʆyK �7�'|LG�7-f����\�����@yRi�wǌQ2;�"a�2����ab�4��o�J�;����G]dr�D�h�o��;-JV\�pi���$�I�
����&�xo����m�#D��Y�Vyfe��ɢ�M��9?�:��"�t�g�b�����t?|̯5��z��{���A�Z��d��5Y��MZE^^6��<���|>zS���)�t���-o]�05Ԥ�"f�wM֍�σ��L��ϧϣ��ͥP�`�Zn�uS{JGAV ��y9���!�����5�'k�=�|^u'z��k%��Σgvd�}��0�VB*������lܛ?	�LZ`E�9(�͆_�Lx��E�4���W x3H+~Z��m9ƒb4#\�/-=�t/�E�w��;��sVM��`����Y�1\yX|�"H�R�^|Mg����yw��J2G����iS0n�h�:�v8�~�h	8�J����`4���Q/qC:�멏�g.��g�e����j�1�1��܃�3b?���?�|Ɍ%ԭ����*�����\,�<Q����Y�/_��A�I��:�����曵-���ß�GN!鶄��,iNl[LE�ůl�B9���E�ѕ#KQ+"�O�� ���3��icqҰ�jč�.-J��=I�G�^�+���i��w���%��8��L��'�~r4��p�x�[='
�����}�ƈL׸%�E�k�~���N�:(�^�rvUe�.�n���8�!N���x�vnD4&x��$-��3��� ��"a��!��ŌI�qĨ��U���PJ8!�:3;dB�e	&�X߄9�~�2I~�#���L��?��ʺ����i,�,�i;dKkg���	7	�De�OA� ���M R�y��¬ш�i#Q[N�rۃ��|w��D��:����W�1~�K��j�:�5�QA
��+��2`��h�F����Fݪ���$��ו3kje$��Q!�[��ub�w�f����Dږ���eZ+R�s��)RX�v|��|1�.qe�Wb*�����~g��ӳ�r�>;�
ag1ckC���pPcrc�|<��$�<7&g�P�����qx+�K����h�c�dHԿ�1[�;����3P��w}��(��yA*�cO:������	h���0o��KC � �g}C�N�<%�U�z���:::P_�{+w�Nu��QS�UU;hl��m�s�fl߾[y�Ճ;�n��m�k�FTTnCu5��U����yj��m�u8�[���TkKv�܈-�֠����'�ڙ�p���zN�*�6\�ge���%!C���_z���4r �ұl�n&q�C��=�!�����v���I`Y����� �=���I��0���L}A�F��qd�f���yK.�F���{�j��ն��~4qO���F`P^�ђ���^�U�ܝJq����_����+v ��T���C�`��"x*�)�F`�7�/�T�H�w_4�4$Z��lh�W���r=�	�/s)Q�|��<�-{Z����.J�����Bg�&w"ܴ��<�5ubOM5bAM$�>K�2c�b��4���Alm8�����C_�w3��j��x���qSi(�O�y��Y6�p��P�7n�%-��B��iG(���f�65!/Ӈ1cGYyXSހ������|1��h�s2+x�1퀾8|����Ĝ[�"�� ӛ�o��������G=����'1K� f�O�GZ��\�����FyOmU�P]Yw��V�9k\z+�
�¥JZbStl���:qv$2��C- f�������@�|����"'�'n��wuу�t���j�$���D��b��X�+����-
ѓ"�مA.4YJ⥥I��YYtɕZ.+�),$sH:�M"Ʋq�`���������k
v�ރ[��^~�=�7��e�f��>x���u��r�;��%G"�/�4���t���Fl���G`����S��S��چF,���R ���F[k#|?5�,ơ5@�*a����\����H8ƶ�e0��&�h����~�I3y:��5�{�4�˩��W���ī|@ف�~|���0n��H��Hк�����ٍ�
.���uk��n��݋0a���3��wc(z����"[[ߌ���z3>_���m��:�����]�Ro&珄7�T�b��|X���$ 4LM��#����D;�k�T}NlK���E���+\'��D����j�xa��P~&z����cG���룑��<��Km]�Y����Rly�
]�a����2ŋ1G���'NGai6׵�'>Ĳŭ�Il�4�%�i�R�x�Z�纾i�F���MM�|��#����k� ��!^L���̯[���|���}1r�)|nzv�	��L�x(Y��t���y����5Û����
��C>Vsi�B��	�v"�<��6$|n����W�2?�*�#<����G&����0g=�bS�s�+O�I��/���j�6�uD��OQ�cǏF<���;�Q�G[Ňm��h ���rj�DB�d�a��>�5� �|>;�bex��!x����C�b��#-C����I`#*���N�uk�@�9ꞩ�rG-2��.�\�+�HUT�.knBG�.�Fq�7��\�Fi$Pl�!��`c�ʗX��#Ļ5G���ˢe��
�͒.ٹ�����9��(���M�]��_{φ��nÊU9A�K'�7ԣ赴6f��F0�I�G
���r���;)>ҍ����#҅��}�;����EBd�!�K}FN{�Ɋ��g�jg��^�P�i���`[ޛ��'��+pF�&�L"�t#*�|In�>?���[���c�i���w��K.���7~��� -��A}��*g���x����z%F����eC���0t��:��=��5��R^�E�(|6�@�g;R�)��(|E(I��������9;�cK3ˈR�������* ��	 {�S���3�?��xgC��u�>^W<��D^�IjCm���d!�Q��~�vƏ��ld�g��`'6wD�tQvR�H˵Q%)�~�d�>�8��R�/�h=}����gi��d�GEK��O����g�2+E�H&��-��8�@�Ӧe�4h]��#&f]�hs��%����-��vSp� ��gQ��Bd��8��h���-L�G�"q�����̄I��H�z��H����6暔3&�(��Dr
7K&����'ޙ�Ê)	�<�o'��љ@���_�Ge���jiY[��X�;	����L(�D8vk��#�M}�#U";��'#�ݓ�?v�J���C1c:��r��Mhj��P����/��H[�x�gx����_��+�=��O�f綨~��Z�^0�R[[��;;�
.�H�Q#����＆�{+^|��]>�v}h����ph��_�os�0�.{�G�"o[:�n�TI���]=���@A~6�H�fg ?'9Y��#;�CN�k�,Z&<�!%�1�ʚ�X�evT֠���Ma�4QU�JZh�^�׵D)�b�絾9�+}[M���iHS[�-|�ڍ�v`7���SM+*h&G*1
R��'q�֠䋒'šM���hTEh�0��h_�i1��`q��4?��ވx�V�Fl�%m���lX]�;��N�����r�cF�xLg��aa;<�1���{mP������O��EY�V�'�����"��7�M��y��y+m��m�`�[5��x�W������ۖ�_�»��Ƕ�k�g�J�_���Yo{�W���<��F|����b��tiXV0�
����Χ.���?�koYKzF0��haeD/�U��8��c)���d��z�[�r���JuF��Nm+(�#1�3����	_C&3V�qȥM.��U��v"P��c�r�ª� �EBǘ��*:Oĳh
g~�oH*�f�~�+z��*B��ξT7f���P�	���d>�2�גh���s�S IS��;��\L9�?s*1�aj	���Rs>|�����O!�y
Ƕ��v�;m�[.�W\�#���7��o���?fh�$ 	�M�A�{v�?܋?��ؽu�i.	�K���������o�{�On�7}�"|��_���� �s����:�[�nE���݆Y�E�"�-�7��H�1>�I#�=ӄ-eB=��%�eF]�,ݝ��9��������m���~-�[�d1�t���%!"$U����޽,zO?M�&�=
�JK1y�Z9�6g�E*i��R5��Z��ܰ��!'fC8܊��Jt6'���$Ļ�E��)ʏ����vF�(5ʢ�	|�:]TC��NLh�J������qW_4	�(g᪳y�3�!_V����*o���
K���ꅲ�!:k �C��j�`������� ���퉘���(����%���Ix��?a(��D{�b���W;T��2�a�L��c�?'��iQ\\K<:�Y��F��ń�(Ѫi&�ƻD�ZC������r���w��5l��`n��Pഡ����Fd{S���EP�rh�-)�^���,&u�쀷�D�$�r��g:���I�����U��J�Z9	�AEo�/q�r%����N�ԑ�Y~z�.A�DT�Ё��J�љ3��#SiBT�ׇ~�rп���h:*�M���Sht";+c98�?�4�t��+�����/q�'�"$�U+��{����/ƞ�6|���&\��x���Ι�'_x��� g�}.N;�\y̱:|�	w��Xo6h��=x���#���������ӑ�&�6�Y��y[׬��'���N>+��Dm}F����^�Ks�2ow������8���1�h+�,��+I�/�S��!+?M��p�9���]�Ia��[����Oz���r���ܬ\���vDJUS[�ע�f��o�}%��.���T�1
g�}.��wq��c��&��s�*��� ;;�y���~ST��8�$�s���ۯ��U\�=�J���L�ܳ��=M5�}"5�O�'l�r	s�T�k뚱�b/�5�D�N� 2�H��F�?C�P(�m[�:݈�kE��ȂI�+�V�:XNte 㪍-����{V^l��<�OL�0,#,�UgNƹG�ñ����3G��YCp��!8i�P�t�`�2kΚ��كq��A�=y N�<�0��3��i�q��1��AW�� -*�W�Q��|���,>�N��	C�Y�Q-�x�q}����n���b̀R��]��l5��.�#}g�m;j;%�`�*XR�^ԙ�Qd��1�=�����%׌񽇂H@H ٮ�	sU�O��J��1��&����drH.�G��� �O�HZUJ'�g��G�
O Fw��	���gu�t_-&������� �"��W�--R�涰�u뎶��m�/�Pҗ�=���d���#|�c"����]��K��'�ޙ���fD����E�Ӗ@��Ze�2O9�,�|�i8������V��Vi�rOz�a<���hhlD�����v�VUC�-Ēk�n�fL�}���e8��30����|�v,\�:?�_����:�Ǔ4�J��ƾ����p���7|��v-�}���9���'5�x9G�����N�d�ޥ���s�[o����ι�r�sq�/s_2�c=�=�c�)]�4~4���U���kq�ga���Rõ>�X�&������3&��O�����n��ƫ1j�0[�ڭUo�?�{k��Ae�[����}V�ڮ���R��u"���a�-�VbӾ�g ���+Lk��8ݛ'��N��F��½���!�i�4-��*F̟!-�M��������*������1y8i|1N���f��!�8yhN��Sp°lU��Czeᨁٌ����px?/��1�>�2$@CE��,S�|2g�몷j�D��K��).�Vuu���5��P'
+�����$N҈CZ��oe����?� 
fi6��m��l2뤖��t���	��ћ�H 壬`�����'��N�8NX��(p,��ľ<�Nڟ*�4�{'�\j\���L�5��N	�Ur�W�$j�|�J�?!�)7�dqu�"j@���}QmG]K �%˳L�ԩ�h���Ի��|ڥ9�*?�ggP�uQ�������U{ym�-hT���@<��+{*��e�V�k�v(�[�z˳}��t폷v��ڳ����!пw&4�쭬Dg�����.�u�[g�kd��>�?A� �����~�N��q�|�<����8��n���O��<\&���֑���mqA #�����c�� �JMf��5����N����y0d� L�:���!7;�|5l�o��S��O�5�þ�EدJ{Qqs�N�*��sn؍ξ�Kq���E�rD�p�Qږ+3+Ӭ�X��4��N��a���vt�1�6¬��O��n���$/��8,��5y#|�������\�#ƛ�����(��~��h��0��ҵ�v��6�c�q|Fz���쀌4b�U;�g���<HI~2�@z��иI��8�w����8y�,���y�3�U� I�d�{¤�3���ϵ��	��w]0��U-ؼ����h����A��Ս�
��zR6���Q�Q�SK��%#������ޑ֥�e$L�%�4k�GJ����Nl�u�[d`�Bɸz���1me��U)	5V��95�&
��&�;7b�d]��y>�6�|!L�6	J�QΖ��T̄�	������m�ay������D���ȹ��A�O�k�KNN&���x��Ŵ��X�hΖ>����v:uM���@�Աv��|ӏ��on����!���%k�@Ar��?���<�s�u�s�X�=Ve��zu�Z��I�"חc�kQa/j'9��[���u.%�?���������y��vM0*-�w�:(1;�on���;��R��0�K\�3�]ixu쀊!��{�~��럾2���ҶB./�zJH�� ��3� ��� /��i�l��'+��.L�g�c&��d����z�-a�./�/��j7r�0�6)aN�ix���H+�<���b��h���y�1���O����Y�Y(((��Y,o��.�#1E��b81�C��7|�w�K���R���x&N���6�|����-xy�&<��
�������>w��b5ޞ��-X��x���x�5x��X�a��ۈ��q,;k����UX�Y��E����܏�:�<qu��@�w��^(�%�e��r��UmX�7��MT�#��bM�P���hUj7�wc�<�H(HiED���@2��mA��B�'IJ�B�Z����(�C6h�N�k�Nd�P2qy�0d�g�ҩ��[�A���b��Zː)X��G^CB�B����p�Wy�jZ��
�`�έ&јya���ck4M3J�#�j���%N�����v�V�fݙ��K�a2ޫ�ښG-�eNQYjf��7��B�u��(�U&h�F8\}�Aee=6��FX��L'6�݌�>�n��X��
�N��b>� s��8�)vH������L�iG�ƣ~y���5��(��Ȕ�lo'�wv�z�׳��WsƄ�zI�C�Itk+��\�;G%�KS����s�a��%�(߂��ݨ�ރ��J�QYq�jR�'��[��X���:4�6���
�{�b��/�r�Ǩݶ�JR?�$����q��0�V�!�ƣ����n�����v�7�a����-ATF�O�-5ظe-�-����%��`��ϱc�:�5g������_۩�Y&ŗx��L0٧� ��;��S���d0��0�M�z3�~X?/
�z�ȟM+B_`���|�P�V_T�S�0I>�� ������v�O�9�Ɯx]�%B�t�|�GĠ�}�[;�P�(o�ß�������O.��O-¥-�w�� ��q1���/p���?����\�˟]�U5Ą��+oK]���Z<��&t�3_Z���݄���U�hS#+���Nq� '���t��k�77_%�Ӓ$�n#�l
E����8y�xqn��f��������%m��]�32��1e"�W��B����4d5��J0a`?e�|T�$,�!��T	�KE�|�^�M�Ur��Q��ĩ��Ŕc$�I.�V#[���6K��4��V>�M�a�fWŴL9:�T_{W!��^U��R��������:��8x����3&�ϡV5��@(��	�uF	�A�/�?�|�<��۸�Ƿ��9���xU�+7���<�2hmf��b-��{,�R�"����`0]N<j�ܸ�K�1p�X�q]]�K�R ݿ�E��;�C�cv7�݆�}N�}ꩧ��߹�Lfµ�\�_]w�t��㯮����	���Gx��w`���Ǔ.%-f2ʍkV��{��=����������/o�}��	�t�Mx�O�`c��ag�o:��,L�x.��ո�����/�����l��#wUaJ�Z�p�V���-]�?|�{8���p������9�<�6�8\~��❧j���|�{��e�D�1O�6�y�W%�Y�nT�p�I�d�Ѩ�Z�aq<BJ@�GzM�-�okAGg�jjPQY����~Da�ݫ���OW�o#+�v5��[k����ϙ��]Y�]QtT��iK-�hXт��5h���֡}N5ꗴ�iY+Z6u���è@����vc�]���n��]��Ga�����<l���������Z��
Ż��ņo�α	�33��Q-�~��"ͦ؇�""�7�Y���dd�b���ɶ�����46�1n�#���
��{gD*a�d�tR� сN�ol?$V*��&ԙ��s�'9��vs�B�sIxTc�$����w����R���Ж7yekk�� �1��wR �J��D�</�������L��Sc����O��d�CU֋�X�,���9���2\���p�)'��#g��3N�3g`���عe�����N��"ÆM��I/�S�0��h_�t	_�njs���V�e���Vy���T}/�9��?��<��}%g���I[P�0E���H����\ �7t�5?ďn�1�������Iy~��m����x�ٷ�??��]v��b9(oM�~��|��{q�/㞇^�=?�?<�"x�=����$s�n�dm�C�H��(
��ǟ�Ï�&f�p<�����i]�#"wI��i�aޢyx}�jl��Am�^TWד�ס��5Uxga%^x��5�D�\��v�A�*.j��t�Juu��+�E����v�4��3�yt"���dү��sU�v���I�6�>�j�T}�
o��Tu�~a��lSks�1�ß���Ԋ'�дr*���#a��d���e+a	� �EA��H*�������Kˆ�u}(�>Y�G�Z��y��i'�.}��4�VF3�?�`F["nw�*����y%�� �U�ו����g¬��ŋG+�b�
��5v�Ål�/&��v�E\߳� m�c�>2ˤ" -?
19+�?�s?gHg|�l�W��I�d:&L�d��җ߂q��!	��wNi���ʛP�5��JX)���(��L@jD�'Ʊ��Y^�'�����fٙH)d#-�F��K�� $�b!Vo��R'��t�~l`�b��G�B�2��-�Eii|��8��()(@Y߾��o@����d�XADM�3�>��7"�RV\V�x�~�AKUjwU�L�5��ko�ݗ��e���	N�[G������;Ѯ�sG IZ�qD�h�����)c��!�9}��ۤ͘��F���vзw����`ײ�=;�X�Y[��� @������1n-���v"�C'��z�φ�t���H�90x(���$;��}�����>������}� �%�c���4(��B����'F/&�b�g��wcO]9��N�#d���r85$Z~�M��N����e�&��|�����S�cjyR� ����i�0������u�����5i��	�~�T���g7Vt�G]p��g��7�ω8.e��Y,��3��W
)�隃� ~�7)��5*㊼z"�JE]����k_F�Y���%=$�	��<���|�������1�򢃈hؼ��`by�ӷ��|%n�j�0ъ�2���[f.�c�WE�E�#���H(jkl<�^ 2�	���Sxr���r�L�uCdNI�I�3�Ԑ��E�S�T\	.	��V��]��_�2qۏp��.B��͹Fp��`Td5�<�ڸ����AS�%�-O��z���~cQ��G�Oy�j��T�W�=��gQ��4.ޫ�:GEpY;,*hih����e�ji�R$E�+bGh�hY�n8�yu��`��nBs]#��%�2EPi����LdG]���x�F5F�[�|���a��������K�G�*��ӣ�0�ka�7��ӫ�Æ�6��v�#eÑ�Y06���|���SZ�[1��񓢤�=�Z4C>����=�eǙ�|�5�O��ɤ��1�:����03=9�y���pb��]�b�v�F-W���B	��I�w������R�Ti����e'3�У�I�(AF�v ���W�6ԯ�%�ا��R���0��Jx�w2RӉ*rL�f�<D���w�O�� ��[��r	���Ӊ��K��8��+���"1��{�Rcl*���Kv>��x+E��J4|&��i����7n��դ}˘��9^\y���Y	:yg
+��l�X7'�Θq�J�0�V��?R�d5�������a�	�;��+}��I�[�|�![�f�*ID$���x�ȅ���6�Z�"f�BCf�!F $�56���07�#��� �$a-�1�'X�Q\��u�qE�UGM
#�����l����*�y�V桟9+����f7�*\H4�&`׳�QZ�CsIQ��ɼS��S�l��T�$�XYK�l8UZ�Nd��N�Jsiu����݄�iE�CM��]�n-����ʫQ�vӅ��T���d�W�2+ӈ_��G(GzNJ������>�JQQ�{*w`o��Y�5u{����4�+���I������vP[ٓ:��#���א��h���8Gq8��>\s��8�����l@���Ag��C���q�Y���^�/��n��ϸ����ֻ�Íw����<`"�U��2bf�=m����z�Ȓ���g�q2�y�9̝?�>��>�(��-N¯�,�F�.G
%{�B�GA�!�(�}�d\s͍�����W݈�ގ6m��r��%[q���;r���©�H��ɼٯux��>�Uˬu ���*d���	��+��A+.��N�����kT�2�Р:��.@}r_�gp����:��C�̪�1��v-L��H(@h M<PB���h�x�?c	�n�r�6���>*��d&��@x�u�Yt7yL�<
�T�#ܮ}�F=N!�d����*�Z��^���?��W�e���ͱ��CTj��K�
���2@�c
@'�q�`�jt5xL����M^e����z9@	��䍘�|r�H�I�I�r7�ZLRYJ�o %$2�U-�W����%�Q�PϏf��"
�H���P]���:£=��w�e�/s�ZV_�s�D�I�Ӗ�9���?���EH�����/��/>���ý��#O�����1��DTu��H��1!nt^�t����3x�`����_y��z;���_��'��q�̙���o��Yt�*������͋�0,ot�>#,�'Y|�$|������7߆sο�o��Ի�"l�(Zi�����4�ׯw1N=���e��W\�^�m����_��x3����8�Ǌ��d�2EOóf����������0��1b�pZF�
��ݎ�Vz
��� �9Ja�A_
�[o��>r/n�����1pp	��pCѪe���Qh⟕L�M���iF���\�m-�!�k:�7��a���#�t�9����<i��/B���ށ��fۑB�i
�����ئ��|��腼�☹0��C���?��@��]<�wd����	 )<���3=���،B`l��ѓ22��,�����؉��L(bR�[.�����z�}e��Py� H&$5�$e0��GЉ�
N� f�G|BLG�h����g�2����@�
���!�N��4�ې��w>+����QY0�2JD7���I��SG0���nU�s�`�Y�,b	�&)d����������E%p��vf M�K�&�Y4�/:�֣���V�i^ː� �*our��1��)�����p;V��DM4D�(x�5�6q��%�8�rV=��2s1��#p��#37τ��bӈ��~p�	g!��<�h�{�5x��0z���L�w_j��/�q#n�j��!8��(`z�jE,�� F��ξ�������>�
�{�L�>��\[&]R���뾲#���7d�T�-8��I�)�Avq��R�A�䀂l
�q8x��A�ӈ�Jb�vDbQ����,Գ���!۟�?�*Y>�]��c�Q�o��,��ef"� ߘ��H���Ĳ�����}t�����٧´̃�N��ȴjS�+>'OC���f�A8<~'��2;�b�����Q��RR��E�5�p�¥�-�YTȼ�)P�)j�o���h��@%���R��J��x������+�[�0a6�͘�����|���S|K������p�H��n_���1�~y�x��'�N��?;��T<��o�_����=���x����g��+N��AQ�r ��%?5����gaĉ}��0�%����tV8�E�j_��M�Hy��+�{(��;���7�,��|#&>���$Hdd�t<>�E�G�G4���uԪ�a"�ϣopE�*�dTB�	�'��5v��M�K$
�I�JcDHB�l5���)PR�y(�K�K'q��GA裠I����[+�B��JW<���	#	M��F¼�b��G"5��!\#3`�b�6�Ma�듙J-*J-$�CXY'��Rk����7=�%N%Id	K
8��I��}��Q�cx"O������O�|�����p�On�?�G�xM>�p
fƕ�-Segg�#fഓO@q�������d~qv '}�������/��^�ݏ=��ߜ��,jV�6��A��*s�$�n����T�?�k��!���:���+��R�0eH��+����.�J�U]R#
��r��|�IEG[YY�K���䙕Gk���'<�a,-���hk�+����v��d�����Ţ�ha�hK3�eh�ବ|�1A"���iB����O�Wy%rv��\U�;�l�"�T�X�dOUn\��-�	�3@�9�ԭ��ֲq���Ά��L'6a�̀?�L����io7O��F��:m���Y�����Is!L�4�"Ru~��F��NB�u�:^�p9�:)�6:dm(d+>y,�5�fP���4L�{��>��ċ�fc��^8��^�`Fo�?� N-�ӊq��ŸpF|wF�;��Ϲ�f␒4Zt�Es��c�-��`Hq:��=	Z�iW���F^�� �Ъ�e�x�0��g��U�}�L(�M/��4�8K�D�F7�v������ƽ7�Xe��[އQ�Vd�۩��*�Bsk[��Y�����u�>9�"�w>�If��f�0�޻%{��O�T�I-���K�:��#1n�D��3눕աu���l��B�&�-h�6D�	f52�u8aP�K�a`�^�߷ �?�tԣ��Yj��6���I�J�!\:�:@p(HE4FX��Β���_t�^�d,.�K9�OC����:3gNǤ	cQR\H\����J)H����Ȥ 1�^���O�=�����	�Gb����[RD-99t���s�����g�����8bT�.�d&�#��u8���V��biR&��?뒸p���+���������r*&N����r�q��UUU��^ya&�O�p�TK�JȢ�N�>��#�;;�w���6.��������^F��߿� \t�q�U�b�ر̑��D:\,�ن��(ߌ�훱y�jlZ��6���=[��|*�mº�K���{~�%��6+q҄�;�P�s7Z����T�P�9��TL3X'�c�=��J�͟�9�HK��P�cB������}Tڻ���p
E��܈��&;jb��rt�Qq�"��R�9(H�D�@暃��0y_B��Ѝ|�hE��D5l8M�&�%R�':�0KǾ`q�S���8�82�`��TF��M��N��=���G�M^�g_b>fd� �}�y��^�h[��Z}�N ��'?4�+U�
�� �A܊��QeJ&HH������T��|t�嗬�9^�6��l�fó_l�u�-BӶV&�&�A. f�ҊI�jwT ��g��Ё�5� ʼ)	�0��2�N��n�L�=x�S<y�1!B'�ͥ�4����M�9G��-��F�4�af��h����1��g����oBg[��*��q#�gcՎ:�쬧�������6�6����3_"Ɨ�YS���CF���ǲ��X׸�(و,�7����3�c�A�KyQD�J�Hx�1���`�(,���T�0�U�c-��D�6gCMP3��4ڍ�F֕Nړұmd	*�nJ��=$Y!r	�*�Lou���2S��n{��g)�F�7�dt!��R��;)\R���H}���Κ����UW]e;�7���z��|K$YD"��/f����_�k/=k�k%��%	#3ۋ�f���G���.����� �5���\���{�>��\g�L�/�K/��8�T8Y��l��iR�X����w��glY�
�ن{��F����$�%7��7�tz*p��>]r	FRA��܋�<�0�{���G�]���*\v�u(*��%���|��W?q�����b��x���P�{+
�2Q�{6P&F�Ҿe�YZ5u5ؾ��.݈��-�6��Hf�/�����Ă��t����ز���B�j����N��U�6zDH���-���F��6�D��h�i�<L��Fj��(��Y�B6�qf>

�q�.�B6�cV ���Gu0��y�?Q
�4�	i�!�X��핸볍�ZB�
*%�f���ZJ��� ��v1���BX%
6���o��ú���]X�uS�u�0��	#�C�bZ��*}�J�I�hK�E-Fs3J�Hd�Ͷ�:�J2��9U.)P��$fL�2D���Nq���t�R�����;��5�
�2���o_�	A���PZۃ�oh�C���r2n��o]:�3;_�Ne�T"�9L�
�IA��H�����L�He~�j�zИ����0]5�Λ4��o�.���#�Q6��^E�AA*��o8g�$@mN(ԫic
W�@�Ome���W$��e.�K-�4,'�N�5JR`n���I��)�&�N�Ƥh�ӣ-|4oFe��H{�uj�?�%��\��D���Icy�3����0Z��U;%x4|,�m*Zۢx��5�����Ɠ� m�q�(饮�.�+ד�/��Mk���ń��Q`۳���<� �i��;��'�����XHe���D�Nͤ&����6l!�VJ%Uᠩ�q���=���:G�xJ���"�vZ��>�gTm�B�Ew*S|u�TUKC�ډ�w�vZl[�T�5�Q��kl�E[g���ojJ�V�� �#�g;k�>��E�Z�0J;��~V!�ǫd�M��r��ٽ���.���t=q�NW>$_[A�'��7l	⩷+pۓ[�?��w~���|.��\��V\��f�{�*�u�
���*���*���8��%8��%8��y��+�����
ֱ��e�I�,����`�Ҏ9��g�#]]�	�R(M�Z|^�O�+�Í�s�^c�Z�Қ���1_b#�G^H�8=)�~���u FB"5)o�%��{v���/�{o{���\��p������������{ŗ�ɅڢD���T����!
F��B�LG6��a�R8���Q_7C��j��@ҙ@�r'���5���IL�0i�V�����^(D�FbC�T�1����qj��a�7AN<j\^��l Y$V�
�B��}��Z�#fg]K�b[wEi�wi���S����K�ʪ�
je�q������6�0��?��=O�����pgB�Vc�c�G�A�����v�{�}hm��կ�s�bK�[�TD�j҄�]�/��H�1��|��>Ck[뫙��6b:��,sћ���hU��!<䢩�o�
��KAN��^>K08�XԖ�]-�4S7��2��S?Ҽˌw��.7�̲��i��-e����p4�����0�&F�#h�A�Ť�S��tѺȅ?3ۆ�54e�/�7�&Og�F�Bĉ�EɆ#�Y\�� �+�Hgqx�{���l1q=�ȇ��\m�!��5��	�J*�c��Ký?9��|&��T<|ݩx�����g����ų7}���-���q�U�'�f�n�"M}��YUyvU���j��2�44�+']��'q#�^�ju�H?|토D��Ϻ�����wo�~�98�sЧO�����dbi-;��L�ۣ�Äi%�cѤ���(~��*6�@Q�J�xz��[�`�W����C��#�s�4�F��aVf ����ɦ�J  ��N#$�tl�p*B�N�*DFڅ�$2;�Ά�ض��Gm5�,##1�Ә�"l~�S�us9�QEca����ՌH�Q�uU"^��۾]_�H2BȪ�ť��b̅�Z�������XV.j��y��wP�}G��c'���I�hW'j*Q^����]aqm��rq�Lg�uu�l��2�auD6�#;�_!����'r/|�.�H�G�&~&��3,����;vn�7��O1s�q7�Aj��@*��S��م��8:�W�ڴV�M�a���&�_�U����0ڊv���ހM�a�{�c�Ud�i�49%MD"?�"�j]�Ai�dڄX��ֵ��v�4�Z��>���?D[]=ߥӊHE:���$3��L�K��U��5�ޙ�S0%0�����_D\�\�J74�W��A�>�\�3�d]�F)4:�E�»��)1�T«�YS\]�)}O�&oW����>�\�w�.@��W�ϖ�1�& ���@D��F%$͟��~t0��0������b\xp.>�~r.=��>0M���c�8y����U'����􋋨��Mwvj����p�d�����	ߛ�{�@ ����>gt��ɼ�9�z˭�ܾjw�[S�PC������L������%H���{�v쭬FG0H�؈�$���u"!�&��\N����ښ c�dgS��+�T�[E�K�9�'���e��3]��4����|�^�>H����B��8���/+u�Z��ƼX.A��C�Ƶ��������21d@�P��h����U��T0� S����É�lK�h&�����e�2��T����KQ]���f�V�yH�j7�	�Khoݺ	󾘋�kנ���5^?5���!<iq�ުJ,���Ο��ݻ�ɲ�ʹ	H5�{)�j[�l�R|��X�v�i���Z���|$s4_ �^�T�W��n=�|�}�]X�|�-I�ۯ?|Zť|�M��q�Z<x��q�g���܍��ʈ�̼<v�T�	�m�op��D=׮Y���z˔-�"��>�0L�1�t���e�R��bZ4o��_AEu]�O��(J��3O?]�C\pɕ�9�d{�N�?@}]>��lٲ�؛��.*
�M�QU��W-ò���h�'X8�s���M|�������cf`�1'�4�-����I��WmK�J�3pġSq�3���%K�r��X�d�����4��0,{8< ����o�Sg
�.ZZb�_���J<�y��!�Z����ǳ�y�l�Y�����U�YY�vRlmC#v��m��@���)d^����x�� �&�Cum��:�#�L�?�'�n$��T�K��m��l�<�;w���*��K/�.�%�k�\Dj�Wo|����ߝ���ß&���蕧}�*�Oj{�㨹Y}~2	��+�������T.�T��(=������ �ۨ	�ʲdmh%RQ�X�6 `�������
��jQ��s�����W����U>M���%��O���� ވ�x+���V�����fL�Y��%�ْ 
�&�%����a�Pő���.7�F�$"),.�7Zc�6"�t{�)Dm�4ڱ6��i���r�է����:��ԑ���Q��6�h�Q�ܻ���E��C]Gvw�al�~(x1(+�&�Cᐡ$f
���'Q������}�v���_��ǂ��C��-d6��C�涸��ņ��q�������%>|��^0�,�������� ��U�x���;o�ӯ��yo�E�e#G"���q�-�ZNs�.�/n�{�I���Gزz-��Ч����i�����Տ�(��G����_í�݉u�ލ;���+��S0j���,�qw�.��~}�	�{�Q�M��,?��Sf�B����ot���ى���@nR�8���9�0L�>�4.���n��G��OO�O�jo����&KK���	�p�m�Ĭ��ƐA���P�Wv[���X�6�6lM( �c*�k0g���|��x>�d>>��KWnFg}�u4���N�>�D�0޾�/߱�H� �N=�[g�'�ޅ�O:�'L$|T��~��ظ;�H,?��&���}��5�������F�P�-C��k8�ZM�������>��S��?}�<@PY��N;��'h����§������JtG�@K�����@>r�YU:�PSBMm�7���F��I�T�"^Mаb�KF/yb7=V��xv���9���G���C����o.����>�ڕ��ݴVwR�V6P��cGUv�4���;jkQU݌��UX�s7oޅEP�B���#���O�.oX:�˄Cf�x�@JF3��,NZ��BL�=�5$�ĺH�	%JhW	�^�(l�3E_�ju�V<�����#�@���Dee��q&4�#Za�Lb�;����'K�\݀d��d�@�eb Q� 5N���8�	� ��Mn�&�U'l,W�:�Z�ZP`P�,S���4�Tig݄;��� b�j����^	x�FB4,ѭ�k(��{���#����q{�faL�@�;�e�>U��1�UGRؗ;ͻ���>��G�z���+�B�W�g~+��7|)����ֻx���ѯo_u�I��=/?�}1�V�������m����h��������|+WlçϿF������R����#�bђ�8�̳���F3߽���c�:��
7��ϰfaNqH�.2�_��kTU�ńQ�q�Ooř�_���B�|��������R�۸u^{�Ӯ~�	����8���q�ko`���F�*.U���h����:/��P!"��(k�T�.wQ�[4��TQ���g`��i�?d���h�5���O0��6��Ne�R�S�ճs�Ӈ�٥9=a$�ꋲ�\�? �'N@�޽���4zH?1}*���B?F.Ä�#�8W����a��p�̃ѻ ��"�7��[}}-�h�1/V�[u%���N�V?J�;)�1l�KGx3�v����$p�O����i�D�-���o�DX{S��Ã*��8����0rmR�f�}ף�ք����h�V�����8��'̈�[��*�"�A����8mB)�|�cݖ����e���p��������<���N���s��8��98��%8��e���m�)�EƲ)���D����-z	p�i@5g��%��@t 'n_Z��?�k��ɚ�D|G� ���eI�Ҵ|�O�	�t�Kv��w&���!�z�lR�ϧ���fb�tj��ju	I�(L�œ��]	hY��K��1��UT_w�T�����y塏0�	�4}u$!��cҜ�ȋŬ0kdUڑ��t�!�0��'zq�%��|�"녠�ӕ�ѶB>�Y�n�܊4��,�@����Q��UOL���?w�;�l]c3��}�q�ƙ~5��~���hn�#Nbh
����cF��5��?��{ΩH����W�@S��檵3�U+WcϦ�8�p�e�ԋ��������%ػg�����I�QWU���>߿��t֩8��oQ(�����W=�8J֎A�7�{[�M��G�7�q'.��8�³p��� ��Ǟ��Ԭc�:*�F���;o�9��u:|:λ�|#��^�:�K���;�k,�	x#+cP�i�j���=��F�
#}��eI�"��h��E��/�j��[�F���,}�G�p�܉�T��Vf � o&����t����R���<��]@2�)�4|&e��K�,�LC?��fM�7h��6D�!�"ZCb@��m�iN�|'�*��|��� ���D�����W�vD�/X��A�-t��� @����~�	���{j��g���5C�G���%�W!N���/��Ra��;��0�je��4A�^W	Cyu >�������<�8�Pl�x�`Ѻ*���x��U�z��U/�!�Y����YM;P��-����9���R�N���V&,�L�PkVJhq8~��$�ĭ�YTc����*�<������sI�"Hcw|�B-L�z���X7[������K��%04/$�֤�,�4�&���Ba�Ӕ���Po�pH $�fӷ<�3�q�@Z�IP �r��8���\���QL���:@B�Z\��������+ng�ȫ\[�C�v�Ֆ�hja�7�:��f։V�H��Oi�����f*wUb��%8nơ�v�A�W�������~B��B�3}Jz���]��_}g]pJz��"�]AT��j���vtb׮�(��g�}6���}з�/��������hT��KK��ňзW)�0�U�=�5wv8�	7�&�����eǌ��_~	7m��'��l��.6�i��ژ���| >��c\~����ε�A�>�kOC-�|N���H���5��ٮtB�N�>�P\�ѻw_� �����p�:��0�V��ȈQ��l]�A��N����׎��UZ��%�Q����L��R�NEȟ��t�1�`��鞴l4�������C�����X�/D���lY��=�4�{�A����x��Q�n��I���%ف��]��c�E��4t��x�M��x���m��E#�1�������ߙ����&f�H�;��hv57aWS��N7�"�����jŲ��.�U�M5c(yU\B��j�2YM�N����K�h�8^�K�{5�σ�)p�y����e(c����U�ËK�ꓻ[�j�m9�#��Rj��n⸎� �G�G��蓙�V72o[ek��s���~�g�;Ǔ����N�8\�洀*ɷ]{rxٗ����S)�$��ɗ��𘬙h�m��hi��*����Z3��Qsk+PUU�k#j�֠���V�I��ש��%��l�U������0J.T�j8-P�؂A�d
7�E�9A��U�!I�W%0탚�BjűWt�R����]�4����.�L�1�Y9(**BN�&�5Y�M���:Y~r������NL��6U�րI�N�����~|,'�[�IG��& ㆏��!�(��X�h.�|�-�oۃGC����ⶭ~�i�srѯ�>�Lğ@��Zl۸:O�04�:p�@
����X&뙟�I��a�Rt8t�:RԃLmǾ�r3���
K��%�bT:�k��ho����e�JՇ���1#�Hl%c�e��a�ǲ-��>�I�������I*Y�*�F�p�!�p�M?��／�y��}�×�wN�5�ez����]�z��qi�ճ�F����5^~�U���38�������#��g"���v{Vij/Q1׽���4�7����]�ؑ|T(��ؾh�L������܌˿}N8�B\w�%X��돖��5�:������%����L%|�q���E�D!jkW��ߛ�IÊ���5?<W^q�9�|L)�H{v��n�݋�v�O�bLJ0'*� ��*�Q�J��(�������y��ZY�W^�:8		JlCO�'�.�I�b�_�����3�-ߊ^��j�#��"'}��,4�o[M�p��.�o#?l_
0-7^��%=h�M�o��n�[Z�Bnj��,��+N�Y��K���5a�O!�S2��E4�'f�UQ�w�coEM�P�]����ʽU���C{{'��Z��҆Nͱ�w �c6֙d�@Y&#��f�KB��	p�61�{V�&����id5��Η[5!ð���{!H�F�Q�#9�e����3Za,�f�>,�6"A���@j�K%�6�PMuC�[��;��;cǬGKS�-��ӫ��]�d�d#��YjYG(��݄�D�4��{���11�4�Հ�C����{�U�y��a�b��t��P�a�����kN^.R��j�Lo��j�C�6|%�����+�>�"U�V��c�܏i�4�iS1n�Hv~���\7�������S�ecʴ����� �������U*�{�Ef����`���8��8Z;kHa�K$�w(�~�&D��{�/m���k����Kss�R6k�L=S&O��1�PTZ���R��d\�:^�-S�Rg;1O��]�a"�Y���J�@u�R���u|�z�KWb���6����Sݝ-�o��yYi�R���N�f��|��0�#'+�����` �����>e��g	"�a�b�,B�az!R�u��s=� ����ZKY�B�>x��PK%AW�(�;�8TB��� �}�J���ShI`�T�i��h/F%fv�B)�R�|���g���ɓu&�`חc]]Z\�I^0���teԤ ���M��=�	:����1�R-��@�^���ٓ�Uvvbib��Cm�mD��Ƹ�x�����ں%��Y��[��	�MH�i!�9,F$�GV����yR󓬓ph6g 'Q�����Cq���R��0��U�yi<a}k�z�T�T\-	��L#��a2t�Iuvt���+׭�pmN55y-�V�D~��4�"|u�LZ*W�w�^b�$e�8$C^"�-M����[�Hg��ԶDN�����+H��D�A"�Ԝ��M�2T�G'�6�%��n��;
�Z`9�9���%�B�#!�W��x�_�t���O���Qh�������C�W[>�hj?�����ǯ��5۷�W\�Q㴇��G�5�ם1&�҄��-����D8㚲D/Z�vs�t����>�v�&����w�f���G���5,�RS�Hs��ZM�f�)f��+J����A��܌4u�`O�.���+Bgk=Z��h��Ŕ@ML��L�2�M���dQ��Wz���.)$�t����"Sc=���Wv�Y�U��4��8i>B�	�o���ѹ��Q_'���ӆM�6�y�:��+YϽhk�c�2�r���2��4�$�D��u��q���W{�'�ˢd�l�3!A��τ�s�8
~��D6��{��X��7���P����q���0�/���>�ٵXJ7�Sy�դE��<-����v��f�#cxb=L��C.���_^z��F���5��鵑+��z/��x�j���^�O��"�����>FRJ�j�����x�$�62�0Ak�0�S(Ennz�*���Q�8�8�6��gL��$�S�.�
c�AY�,_�@`s΀V�W'n�q^'����GƵ�Y���ڽ�a����m�U�3EK��h&���1?��B�F�� X���\绶p���Ը�L���,;�� �K�%NE�QH ��jʊb8�e������/�,�����cO8x�~���;���և�|�fB�:�喊�a0Bm�N�X|�L�VG|2��@����Rt�mZ���A{�1�4��mu�[k�eNwnh�Qc�V��eK�;Je����c�G!��H2���
��o��W^�/~�L<�_y9����R#g�h�an�$#��$�Ⱥּi����X�t>y�]쩨D��s�?��L�����X��#D��
��/�'/<�5��"?+%%dVYX�����6͟���%�Ce��:H�4��_��X��X��,��>�.���yP_�♎4�mYZR4��է�N�JBɖ�df�Wq1至O=�0OE����q~]gL�����tٟ4���-�k8���&���A->΢]쨈�����G_â�>�O����!�I�'܉Z@Yq�r���N*�#��;�>��z/�tcaJCo����ĂH	� -Ҍ�h��歺H@h�`m�c�&<��&<���W��.)8px��0��i<s�*C��b��(F�<�R��^�sp�>���GI�D�X H��6N��i��7	�n��K�v�ۦ2�5��O��R� "��	�)���glz�]3(2���M�}تf��\��;��A�J�7��X�F~Q��������㿉+��W\v9�u�8��o`���֋$t�uގ�l��t�WD�:�C+����-�&�'�	�!�O� ����
S<�TQ�Qv� ��X{jx@H��;N_�33C�>"�`Y��h��l���F �PV��E�3+Y��K㋙���c��5UN�J�utڶғ|�2)Ն}��P(<
�s0~�X��c0y�T4W�a����V�y�-����$�6-���PZ4}�4�Yw�Jʤ ���h�o�����h�L�+5�Ϻ��\{Pk��gUE:b5¬p]^����"V�ً�fLé�:E�6̠e����)������������g� >}uqE&�Ҍ�S��ݿu.�����{���҆���ݸ��w�����)�eW\�y�=�)���Y	,����g�?�	���v<��Б���N=?��N\|������=�ƃ��o?�*w���_���QW�g�.�3�<��{�}�*�Io���9��l�~ͥd��!͟ض�/�ر{��|-��x⑿����JTi���ԯ�^���PiJ#I���tO��2����5,�!~}p�P��������uؼ���R ��B�4�y�������wI�cF�'TI{O����X �k���UOA��2Sc>M�J��ɾ�vH���{]L ��vnnǓ����OV`Gu3�1��ǯΞ�{8�����ͳg��gO�m���_>u:�����ý����|w��\��#��^��G)$�˻���gx� �T�)��F�&)�i�R8FiIj�Kt�仪�Ѹ��w.fd���.����?%���%ք�H ���A0`����3���8
��z�:bz�~�����h�\�زմ\	?	Ps�2����O0|�����GX��Q�@����4v��ǫA4�IdH����&W��ƣ�%5b���]�f�,-��V��!Q�ztWi� ��\��+��FK_�-4y�2��0,!� Hbi�G#Ӻ	;��K�J��^�^�hZZj$��A�Z��fS�e�j����܊��	�	�<����������	a��!��r�	i����Qb�8JOEa����W�
Q��v���M�l�-4mii���:�2��Lmo}J��n��))����u�w��3/�d�߽�G6bt���k���k��SO`��r���ā�8@��h���?A�$;g���3�l�Hgsb8�)a��,��~u��^��އl�T̜v.<�"̞=#����Nk��,�6l،?��>��λ����P��0z�(\q���j�����G�ª�M�h�B447�����Ӌ�&-I'�Ǣ�aǲ�����r�N�,K�M,F�
~��K�3�ц�|�����k��w�]�-�<���z����}G1�n���"�gHCk��'��i�ef�6��S���5�Q�85���dD!yސ^�0�l(Fe#7����� _Hc�ğ�7�rU�<q�.
d��i[�IAﲺ��N�G6*��F�֏G�7��-�ft��ܪ�ܠ2�]��p�'����m�hl��֍1��8jX ���s�� @忹�z�Y�q��b�q@Ne�������p�1Cq��9��d��R54�s��Q�?)���x��peI���o'P�d���e�"	#鄗|��?	>k�A�Es06�o =#��T�i��̲=���Q�c�m^�e˖�W_�C�>��~/��
�����R#O�i�4�3[c�Ըm苈�I���Z�@	B���MSpS֏,�$swCu�%����,)��<쎑M�T[{����x��x�(��k�;P�v龴�Yc���D���l6F�o�Y4�75+H�ܗ9Ea��+(DZF&^��clڰ����#A�oZ�>��l]��w/^~�%<��_a������7m5u��䠨_?��~;�gԨ1��2�r�TWW BaQ2�7���yS��@Mk֮݌�ݻ��P���##���^�=���C�����Q���׭[�{�x?jkjq�I�@Z2A
�N�KJu����K���7�Aaj*�(Ek[#Z���J13�O�����Bg����	H���������t��mļ��FZ:�Q�9�p��X
�s�G���*�k����f}vf9���8ˇ���c����F+ۮ�5�a9��� T߆T�$Sc�>2km���%;�c	��T2%rY����W^��iI��TT3�ƍ�!_-T��gu̄-.�o����):2!e�h�C��rh!hnG��ڳ����uOFJ�������ɧ�T�Z*PW�i���e"ן������qZ�6��� Ym��;[�Dg#(ƣ�z�<�Ae�����,d�����2�7Sm�<��Δ?�����ރ��c}�x#^�t*��e�!�	�(��N�Ú��4W!�
�a퓅1}��^,�#�M���O\�I�hTϼ��^%���M�k��NWgݛ3�V��� �M��r�m�o�Y��l�L`�j�����ȥ�9"�O�چ��=(�^�k��PSS���5dt4%X(�R�k�G������<����m�<kϢl�1ɹȎH�T97Q�K ����ztDN��Ff&M�1�yIc���4g�o�bQw���K��2��$�RKXmIn;^�J���+��!%f��m�Ė�-�Q�\�Ї�x��!(6�'���в!��v��A�x2PYQ���V�K���ڀ��a���8�G?��'3�n�t���9���_�E�&AY�y���g}��Ç���BY/2!��I+r���X�b)r2<h����ukP֧�6��@�B�K�g���l������_��~}���s�A
4N���0I6������i���ylB;i"1��cw9�n߁��Bةd�.Z� ��������ϙ�(/'-�D�^�dw���f���mۆ�^z�&�m�3�吁E=v���h�z�%�X��8JE^n.�>8���0�V��B��V�V���а,[���6�@V&ƍ��˾�C9iĵ��*���r�bTRyhkjF��-���E�F?�4D]DP�����<�PYjko�޽uv|�4���I[3g�_Ҡ�'�aw�׭c�j��2ha1 �i����3-KS������_�o�'N��G
f
�j*�v�+hjLANiR}9�RK�����AI����ACc����u�$?���ؼu3j�ЂB�0{}'��>��>�EG����=x��~؊0������J�4��
�4^�cS�@�'Q������)�B�d���Ө6
��v�_��:���ha��oAym#�뛱��{��P��AEDaM��aŮ
,Z[�������H��������_�,�f����z��Rw�a&�Հ3k���Ƃ�SW���^�~�0��[o�}��*|�p3�&���&qz�7S��F�B��f/n$��ffc$�����H�"�T2xM@j���j��*}i�\okkg��3� $�J�pн ����M^���q��#�4k�V�J㐥��4<��H�cI��i�IG���j�LW��,�"Y䠬o1�h3R6j:[Q�Z�|�!�މ����1#Q2b�����ǌ���1��\�m��bZ)�W��Ə�!�ڎ�g���N<�\�B�E] �h�����u���+o`��-2b(.��BL�2͆8��������b�%X�x*�/EQ^q��?�^��{*-���<�W�aޜ�X�h5�Ҽ8�[c�a�ڷ?k�ΞE�dn۷�㑇���&C,"�a��X0o��_���>}P����>��͛�Af��W��[w`��%X�`17	��6MHƮ�B�?�m߾/���	iCZ�������n��|��x����UT��F����%�\��Sg C�|���b�F���yy��0�R(����Ƿ.<&B+��َ�H{v����?�ޚD����-3?�&MĤ�F��}�S�O&�:j׭�T8)X;�+�N4�~(���o0H����G���H')�vh��%��;6b���X�zB�(*.%�IW�V�࿯��*&�Y�6�üמGSP2��d�1Z���@���^�\ssZ��0���bc^�nE��xZ;^�Y�7��ڞx*�q:b��&T@�@�`���S���$	}��X�@��Ќ#��h���\�lĺ3,̜YVJϸZ��i�<�i]4��Sw����_�ډn�ǋw��%��&��O���g�����;�Ѽ
ޗ�%���5���:U���b��U�E�z��j��h����](�xo�\VG�|���U�U'�����Ż���J����a ���TZ������q��>t/6�^B�u;�[����E�C+P��4��M�,�GV���Ɗ;�b�P�0xTA	�5�	:�Η&"�%�ֽz҈�[F�����X�v$hnl$q5�tVn>�2󩱤��Z�����YϮP���Z�H'��v�hs�!���`c�N��X��`�룘Ύ��3Nư��ão't:\Z����l��YY55d}{�� _|���;��xȁ(-�giS�����1o�R���;ؾi#�0G�rƏV6�S#��f���U�X2w)6�X�N��Î����!�6�%�",����ΝUظ~��A�3�G�D��c��G�=�މ�*��l�j2�:�,���K
b(+,�3!-dQkL��k�m�F�"H�U)�4ڮN�L������)U�����p�i��Z���L���.驢[ʜ�\|>.���o �h�Ha��R��!��#��jJa�㓧�L1o�Y[��i���#�����b�z�(&��v�18��WQ0�aێ͘���X��m��GSS7CT�YH�5S
��}n��L�:�O
t���]�8��k�&����ߍ-�6��X�&O�/��g��@����.�Ws�V��B�ރ0��w^½�^���a3F!���m�#�O;t��.߃��ذq3�nA�� ��T�v�.%��~~f��'�T���z*C�(o�Em��n�avY��WX?;z�^ˬu ��)�.�8�e:;L����3"�4
M��*ī�4�����SHd��,���p�N�y%��ȳ�M�vH������Y�[�B��L���h ߋշYy�y]�ʑ��b�����bm�?�ŵ����1H�$;��B���6�҂xs+ߓ�Ph�É�@R�K������Ki�R�|�7=�)Z�1��^�5��zyc8y@	����נ�|'�jJJ��E���$��f�Zu ��jfҠ���=	���(�`l_4^eg$���Y�!�8t�;c�&pxKM�[d$�I.w����3�C+-��
}��#L)�4�����aJ��<^c��b2i^#E{h���p�S�������X�{�;�I�|֠����1��D4;yă�4�M��A��Մ��NCRb�����qdj�s����DYH��L�$!�ު@cd$��$~���V$|�
�fTb�8�6�I�5]��p$�p�Pa�|� �Y�,���Oϳ�TGz7G��.����^�J��ձ<���M�p��pn�@y%�&K���>��#�r�)F�Z8�N����W���20�3r�����ēNa
���jm����$L���.�Kw$��m���k"�v�>�|�9~v�X�r������p�����g��ZZ������x���P���d��Tj���'���o�c:���7�PM�p��5���?Ē%�\�~����_��㎇;����WuF�,�2'Mu�)|�z�]�D��t -��2[v}��I�8� S�+�T`ǮJlڼ��Q�BcS
6U� D�/���>d������5�KP�R�=�Z@���zI����E-ʟ��7���e���@k������6s��2��O�^g����x4��oY>�ņg7�sG#�T}[Ōi�j@�<z4�U��~gÙ��Q�㙹۰��#/ ���|��x�� \&|�u�[������̳�z>-j9"��Z�$A$�l�p�T}_u���Ƣj4cJ��q 2.J
h�W}p��.؎��P�E2�²ݪ�ϛ���jdȥ�`��:u8���#s�og�<5Q�y ��J�q{g�X�3U}�&m�)��)h4��]���=-6
C��zA��P8D����J,�Q<+C�2�(�>��S���ySk !ԑ9T����(q"Ļ������t�~�#<f�������CA��4T���ǙdD"Z�F9��Id��8YY�V=�Q�NԆN��IOCifr�1��Oc�����yӧf�!;��lh1?��&��[K�-<��<�'��P)���r�z�PMx�&+�e{�Y�����=�Ǳ[��h#�CԠቢ�|8�O.�}ge��	�G�c"�"F���Hx��)G��l)2��\����&F�SV�'F��FcZ�҉&Z��E[�G�qEm��$��hBe��P��.�1Rлw)���mߔj��UJ�=��_�}mge�'�'�����d�^��t� ��m��7G���ٱ6^_Y�>��� /;^}(M��g%��m�٩m�M�ed��9Igp0H��m`�Q����$z�l���@7��'�2�0��%V��Tq@/|��Q��1�뜩�y�8xek�r�ֆpݙq�eQ��0}�n�w`?|��I��Q�������"kH&<���a�/�*V?�h�&*`N<`�gVI��{4G˲m��uM7���[�dZ>Y��gw��2�vm6�T4QP{��$t5-�hlluL����>���	���C�ļ�m���қ�!����܋Ƶe�h���׉� Z�`�4P�&��|���T�?v$k4v�<b�ٮ,O�KK����Sb��e�"6M�*���kdeKB�UF�c� �[����A��Qd
I����X���Pg� W-�ϝ�R�WMDz�y���.�� `L��P�
F;��qI''���K�=����^c� �PZ���PQ&P��`�pܤ���+�["�u�|'��9���ģ�Eu:�ev��b��*�+-�3\���Բ���8),I�?��w�du\�<=%^����酮�K�1�X"�K��o]�\�J:�I��Z�)���è�p���_�����#}j���:4��E��=���@M���h��F;%9S4Hj�Tє�23xH?~�lL�2#FO�'7�6�����`�X��gصf5r�3qƏ���"����&'`_թ�F���p���Miq	�;�v�,�?	������}ǎB7�ŗ����<֯���~Na���5O-�S��k7�R�}K��b���i<Ƨ�d:Z���)D�̍���O� �{�T�B�H'?�tگ�����Ĉ����\�0�
@�K�>"�C}��ֺb�Q*����}D�2up~|�$L��D�ϥ0Pct15��ѥ3~�y�C:	5!kCo��؉�p�a�Y�Н�4����T+w�'Ź�$���O:��ّ�qs�I��z)*�`>QG�ɜua9:5[����v��+�ᒝwj� �p˄��d/bԴh+�Mh&qw�t�-H��!.J�����FL�C�P�B�©=؁vZ:�%�#b�2~4f!
��p��X���QpI�in��� �񙿄��T�D�%u��6�4�CX�^��!�,S�B��^Lc�B��%6�}��|��-Q@:=Æ�bȠ��Wڞ�ZԶ����\�}P���#��` �Q�:������g�e5���s�)R�5��_S>�X���\Q��4�pPF����c A�j��u�;��-�-:��U5͹�ӹ�Ѡ�{��ƞ-�y0?�M����$�8L^]'���U\O�z���}�ε��O���s�]�*�.	�/��v�ޅ����m����Y$��C����m�I�SV�2�F$�ư}�Z�y�Y,�d>�/�˗,�⥋�l�l\�
��z��;id���6�����Бc0}�L�?��LT��ĺ%���5�>���#�<��w>&||�	{�V��C��������3ѷ� f��_�`��H�U]EE�1|�h�<��y�i�u�1�Ѵ�R��/q�/ӻ>B%������k��KKiy����DqioZ���&46����M;*��B��{k[Q�D$(�ņ�i��Ş���,�ᧂ��T>�ic�>��K��a03�׽�6񽺳��Ęs��a$'4��ŌJ1mL)^���������T�d��ہ����Ď`]F�Tt���O��������(����Ú�f4nie��nvU:�}ma%�QQM��8a��+˛|��#��鶺�+󖕵�*�/S$�So��Y_^�nC���p�V�v��� 2"Adt����{vTR�t�%G���Bu�a�¨���L��6�����f�~����B%�v����D��(��nk��,��onif��h�v"��ٲ���NA��+ϖ���N��N!
E����>� ���
7�M�Xi-��/,E��H��3�}�O�(|H����à�}lح�����ȣlʥp�[��C� ��ǣ<�g��	&�%��@��6
e*�FID�;	Q�`M�HCe�5!T��YR��k������O<^���; u{�;�Vv�w���}Y��2��YZ���G��8�	��b~VU\!|֝��v��k�a^�I����|��8����ם;w�瞷E2�1u#;+?��F\pѷq��CPRR�ʣ���v��>�''�zw��[��_,�_�ϾX��!T�c:%����L�����夵f�(%c*����fݒ��ݏ�t�N4U�b���8�;�Ŕ�3Pܫ7ک%oٺ{+��[z�⠩S1p�0ӊ��Q�J���L/,��P֧�����%����Ry��2�2�u�
���.�K�J��ϒ�AAa!
�����4��|���}�|��i!1NU3�;�yQ��m��c�>1Z��\Ç�� ڻ��3Lj8�U� ixϟ��t�ֱ�z�gm A%&�d���0�DX>B��)8pbo2����z��(/�Q\��Ȳ<줅S���ƈ�v.���O�1Q��n�R>�4e���W��e��ưp�n�C�� �$]��ْiG֎|����2�!�)�:��\�hur��Z���/#����Kƒ����H�U�p�>*#R�|�gEZ")$�4�u�
�/���~��c ����Bk�Ύ.
�(B;;T��I�@gf破�/�ȶx�Px��t��Z��:v�uڰ��j�"3�Q���*�ͭ��k@em��U��k��Me�xt8	���uu�������J��#bKJ��[���kYz��� ��/%��M�}��'|4�)�ө)��^_E7��h؅��=��!!i������_�y0�����mΜ�}�E B0��&6���ǟ�$�6 ��&��͗ر�8n`�L/!�^GM��r���{o�y��ޣ���/������Y��V}�[W�v������8��Nڄ����F��� �����w��wφ׿�U ��y�5�l��u��TRC��ԅ�p��xW��{�B�'x^�=���
��wLGI�./ ��w��{im�1��б�}�z�>��sB���8��\vʃim�ᆫ�Ş=�iZ㑰~M���y�ϻ�e�y
-�L�N�$��&8��ӳ��,�cֵ���4���(]��	x����fY�g��h�`����)���3A�A��[ZZBK�H��'u�9�x�۩'�,�����������nz �ӖS)�t�2�Y��zݺ�l����kR]�^�ޝH���S1���(��+�#u�v����ۯ[]y�{����٤$1c�p��]�4�>�	��fy�� 2����!�̲�ܡ��S���:E�^;��G�t5^���#�3�<ٞ��j�Z'J���5����\��`{�;�<��	1���h�A��U'�Л$'�Z=͚��1��8��Z��̙ucW�X��;k��X/{�?��><����1�d���x��؍*��ꍠ�3WƲ��x�����~�_��~�C���o���U�%�]X�t2�7���x���4���wb�����N���t���Q��o}��p��Ոk@�*B���[_����x�n�-�@��v�8�B[�(t�~	�������� �=:��L��:j�P�C6����7ZJ���F��Y�QC*�D>��0��˴����Yŝ+_I�p�,�e������/��L��<)d�D�)��E6�MՐ���8��wq�Z�B)^Š��a�HNP�c�nBR���-we��`��ݕ��^���N������W:���o���oT}���@���Q:�����Y>'�����y��Wi�gh�S��_�&�
6�fq���q��SOB�k��dd&mu�k!qO���%TK�+*�9T���ׁ�5���g��M���Ïc��
1�"�ʔ��u�\:�K3g1}�8.�}�̪}��"N{��OR!\C��4�T<�_��'oЯ�\(��T�f��/H��h�̩�g92T6�LM��u~���>j"�#���l��ro�K� ���A�܅��S�O�/�1qM��vXUZ5m'�������+M��WZg���*���/b�Іe� r������q�Hν�� �f�/_����rX��"��q�}����½=J!!��6l2�
�e|���S���dź�T;4�!:�
 �YF�y4��:��p�B��Y8��L��ZP<��
�u.��v�J����qǩ�|��sv1 �Q ��賍"Z����#��l12��a�ί ?�ޟ�uW�7A������̠�����_q#>~Ǉq�mo��{m0|anѶe��"�`lx�~���}�{���z��I,--bnn���"3M 	�[_���/��W߂�۴��+���ͺ�/�4i(����d�%d�DJ����|�&�u��J��$LX���G�{ۤM_�f���!x��0[�i\��j�m=�|d-i�N�^�{R�_ة�D�fO��K��t�fiqgO�#w�y�~��}�	,/�#�կ�܈�:%��ۤ=���>��^��SG�Vj�\B.����
��Qέ��*f���4�u���/(z�/��'L䮼~��?+�┋�t���W�i5'?�a7 �'�Ӎ�w���Z��{߻{!��N�M_����ç�Aٚ����rV�呡%?77��'q��1<����_��?g�Q7�&��^�&X*$���A�ɭb����0�x�8�ϝ���S��9���O��}��/|���]8s��(�&u¬�w�Q��1�Q��{��%���y�w���g��|�s-������3�����œGq�'0}�V�g���h�zt���{�����-�t�8?�%T�.��H�s�`td�~�����ay-c`z�uoل��I(lfV瑩�S.0M�6�f�jAu�Me�C�t��L��T�O��t鷘�D��gc���V^��}�W5�$��q�5x��!�C>̗��=O���*-�R4G�^l����@�3`�BE��W���5���j��(�H�'f3��=g�)�$a�F�����N����.���1-�� Ҹ���$Č݊NՕHc�k�pVq��������|��Ө���(t4�\'k�3�L-�6n�\�6}�T"D�8"6�}o--�m4k������YLO/2U\��z1������x�[ވP�����Ξ��3g1?C�"b#(���ǻ�ݸ�Ɨ!�ڹA�����6}������co{^�06�	:�say�.�F?���{wR�W"�%�<}�}��]� �N-���M�g��0��1��;���A\\_�ӳ�٤�D���}	"���7yqEG�d̃�b}�ݒ��sJ$Nζ0m�����x������|w~����?�o~�<��c8�أ8z�1�:y�u�����N�S�a]��JS�cI��ch�Jd�P�=q�(�s׷q�]��=w��<��c8r���9e��Ǣ�3��3��Ε����E\/^O��ى�R=��\O0����Y�t-i�ᔓ���q(ozu�i��*-�-	-�К��sJ�s�2?�핮W��,�����g��Sdh52a��K%�����:q��|
�x?�����x���#��a����j�Ri��J�ws+�;G��Ï>����}�a<z�C�>�CO��|�7����=�K�xԺW��Q+cm~�O�ƙ#�pvz���UN[�nh[�������8��x䁇� q���܍���/{�A<����=���#h�غob�>��n�?�cf�g��G>�r��%B!�
���6T��KC�a��Y������#'��e4���3�K�5����Eh6�/���L ��!�:RZ��p�u1��.k⸞��<+�V�0r��,i�Q:�F%��Bm
��#�}X.6��u�=6K��f�4� F�"�❥�	\X�gȫ)�a�~y�+va8���Y×�=h��ˡ��m<��jy��cx���к�.��ʢӄ�[�*���h�!8V7Tz�<T���x~����|_�*��	���`Y
�
Z��D֮lyJ��}����]���!�I��92�V�E��̨N9���)?^s�M��K�a �j�s�8;�s�Xy9j*�x�u��ַ�(RCc���qaz�D�b^�Hӱ#Cx-��W_c��L��܅�X�?�xX�"��4�����*%6�{
��������Q�M�6�#|��H�g����`ϖQ�"�d����,�<�9`�`/��U��`q��KL��-BP��S�1��U��x�I|���>����_�*N���R�)%%�� #�]����8z�i�Q��g
�ӈ�)��{�R�ʽ(+��hz�2��/����7�Wv_å�y��/ֲ5�9w	O~��8}�8顉d*�h,n�gا���ߋ�O��޻j-X>�C0�=��ag�Y�^/���8Aܩ���4�Z�����+D@5Z��x�{q����3OBau�����?l{�9��sb2W>?�9��т��(��4��'��J�G�3�2�Ս2�g�p��4N��������
�����Լ1/-�d�JW��Z'��
f�6p�qgVH{K\�?����3��K���Q�ӛ(�r6�N���)T��)c�VN�YHyҟ��z)��:f�j�-�y�a9�K�e,�cL|>��L�1���j����կ��f���u���J��>����������"dНN��-���[�`8�O��>��,��]ˠ\.VK���ڙWڔ5,���z§���aT�5�8�u�:^4�g�z����j�^���V�A��1^��7��+��!N������=�K�Z��ls�<�ȳb��%�Q�^=�Eҕx����w_��v��#���S���cs�hs�^������̗�p[z�#�9�<�`w�ӮR�Li��f�(�	 �ѩK�ⷖ��g"�
�~Q-�v���DT����V����L�K� ��92�j��Nq!O�)-A������to�T\����kk���L��	���مf�S/�V$�Vh�g���Gi����L�dEm�\XC��N&�j��E7-�Ejo'�9�l�e���פ	ՙ^{^y(\�:�<��[�z� 5		 z-��i0Rp��J���X�&"hYI�T��R��>�D��^N(��b�'Ϝ����#�����᜺!�k�?�o�j� �B��3����7��'�'�=�b%ϼZڪ��ҒW��6~��翀����Ox��I��7���Ϳ������ݿ�����ÿ�{���ă�������p��)��)���N֔�YfV���g�;�;�;~c3�3���?I��R��%j�PW���|�igSZ�q.�P�:�Eб��mI�7����^膏Z�����g�����O}
Kd:�w�G
�GK�̧>�;~�#�������_�G�������x��P/S-�g�6%���j9��:����ӵ��TA{���)=7�:���oZ�M��1�guf\�ZL��Q|m�8A��'����;^�&����B�8ݐrNe,ds��s��<���Zk�z�-Σ����&Z���Y�{���妵z��M�~L��K�/����
����<��(,Q�]ϡ^�q����<�	rƐ�R�y�u�N����r͍0�u�{A�k��)Y�)��h���}������GcB��팙i,41��Oݻ�?��!<r�"�&���x����_5~��Çy}�u�H0z����'f���N�ba�r�n&t�Y�w�eeR��cT_Y8ݟ�����s����>�K�݄��������]F8l�?fj
��1J3�;�~��)�pnn3'N���3�>y
k0
$�dy(m�w��9<u�0N<��<�85ʋ�S��w+"��JS�~��?��'cm�Qδ9ሦ,JK>Efy��1L�>���h�Jd̴"έ��3籸���5�M�(\e��5�#��ڶ�n"��m���S#�fQ���:�S�&+,����z�L[���V��4z#/�� �� p��YZ�����xJ�_�ة1�v>�S�&��Qs��g��/����ءCd�ek�+�~7g���������������_�E��{۶PI�F|�)�ΞB�Z�~�M�Տ�6\�J<��!|�K_����(P��2Z�U9kQ�܁J�@Fv�x��{}�?O��'v���שD����@�7�A��c�����H���B1��6;H�-w'?u�f�Fߨ�i&�C��'��3����K���oQ�҉�N�����A|�o�g��7��x����	<r��o��?m]�����{��Q���|Z"�C�/��K�r���)�����݋�s*���������s�v_:�W0��7��֞�މ����xt����R�w �w"�Sb�^��۱���%��:��Tb]6�8oK/�)�i�0�s�(HGXkMa#O*VQ�fP�i="���G��9�Gk������.�`��B�r}�.���u`E�a���!a�&�Z���%r2[�f�i��z�4�M>ZkJ)m�w�H'M�2y�6=[�X��>xGN/�ƺ�[�m� >��x�5}
�Q�W��i��{��SO��`v�,;�C��l��
j��?�d�9=;�[���~3�wz/�l
�Yͩ"����P��4x�; HP1`(v�_i֗��:��!mcԱYmL/�㙳�8~₍�dV7l�7��5S�v87w	G�Ǳg�왳X^^B�$}J����g�����YA'�e�l�W�f]��r���8�p���12�K�(f��T(4�㏣��PS� � �I��IFBD���,5� g���ȩWE�A�x��jh=Q>,�1��h�q��Y>"��
�Ջ8�P`~�����/~��Ԝ���L�uq���T���נ�qu�}�+�^���K���Z��#s-W��C�s�I����ϼ�Vϫ�����}�9��~:~�[�>z�6����i\����c'��C���)�F����V�n	����A�l91Z�N+���1z����e|�3_"�L�b�BN\��<�����X\cL��u@���3#�o^
�Aea�:e`�|�_�Z���Y,g�p��y<���X��s.�q�?�[�����_��~�����׸���G����"�PbG�[���eX��\w��K◎��lj�W]����?J���Ұi�S{��C�	��mSJ�9�x����`rt�oކ�M[05�۷�Į]{�k��ٱ{v�]v�؃��vard�@�9(=�=�ly�	+�;�ľ}{񆷽�[��Lx������]Z��0^��]���V�J��RҦŨ^ m;�	S�ؐؗ��V�Hx��#��k��󵺞���쟧�]�?�"��W�o�U�~� 
�@�b<k>;�_��e��"����z��1����n�SLG�+G>��s|q�1;��r�l�#|���b��"�<��?�����P`�A�[y:�3�γ��dx��|kNU02�UE�z�t�{��BI��	B��p���lw���Y����gsp�Ș��8D?c��C�Pd�|W&�n�l�[�x߫�З��|�B+Y���!Z6Y��B���5����t"�I�j������'�Pb�|0�ރ�05�	��u���|�㘟��z��B����݀x"Hs����ags5�r!����=H$0O�h��?֏@4W0���"�5�x�y�����;u�Ȑ
�n݃���Z��x���O�(n,���;�}3����൯5�e�k��(��^��e�/����a|�?m�#橍=��bA������PRL/0�R:jM�v�5W���M�r���Z�vƗ/ँ�;?�����~�p�[߆���C(9�z�!$�I\w�H�S�(��Ïۦ��y��11�	��L�3�_Qϯ���կb���fYʉx����b�.�N�g��	�����{�ˈ�b��|�xǛnE�m�����ѷcxl�D�W��g���_�_���`׵�����E-��`xx��SDb�H�V.#�J"K�{�Zo�X�D�y��.�<s������'X�6����~�7q�K_nuy��Q��G>�����o�^C��PeYϝ��cOǞ�۰�^g�;�ʶ#y�;�����7���|_���dZk׮#��8�k���l����β����`4���Չ�d�^�~2O??��Sy�d�m2^Y�ښE�Y�t<�������)���]�(f�͈pjFY.�������Mі�aN���C��2�������$o�*��նW���9��˶��U<��W�'�Q����m��o
�� -�k�y�v�bgqq'O�M�cr��/��Q:8���4�Ȧ���_4^Z'>m�_�Qm����G�5@v�de����ƴYo�B���O�n�����4��y�[S
0�H8KT9���63,�-	�z�(&��82���<���Yr�Ϧ�T�=�}x�u���=Z �f�ZBM�)��>��/<|�9Y",L�y��YX�t�ru�Bmb���M�;	$YI,�]!\������i5��L�XZ��
6�#�ń�[��1�N�Z����GN�C�6.�� S���>�G���O��tiP�jp����'�q�jS%dק��2V�V��SO#�Q0d�����KQD'�F��uՊN�$�4���V����:Z����A���cfi�>~+s�ڨY;H�R�̶�����,HA���h��r�/^D�H�H�`���&u�p
�P�qXq58���F5�OSw(�\�(~��;�W_o�K���䡏��
o��Ɲo�_w��ӑ�V�'@�@BA��;��vl�Ɲ��/��}XXW��w�����D�H�4i��BQӟmAM|7���+��F�W����x�{ߍ������m  ��IDAT��%b	[͠��?~2+����+��������T����B�v5D��cvn�$��<��i��|���������{q���H��`k����#ā�e�>p��a��l<z��H�@�y�MJ~�k	������O��3K��?�Flٻãۍh?|�y���_�~ G�x_��OS�dpp�v|�-�L�|va�N=���8&v^�3ٵu�țތ���V�5�x��G�G��dNc�/M�~;~��n�B	'q�w������`������?�-dT��ؚf�eKU;n<�q�$&��O��:�؄M��W5�#H��\�n�;Ƭ�Q�/R�P�ZL
N��%ᒾ����O��0}m��-��p:4Niɋ!;� a�]�'��`/ؤzVZv6V�`#>iA�xoZ��3�O���drD�*�d )@ֿ�Q����l�O�R���vEO<v'��co�F�ۂTF��	���ۋ�-;l�Vp?q��>}��A���"��a/��S�:4�p��Z��.��F3�Z�>���6A��߀��+"eX'W��+*f�* �&�;�/l[���e)h����8�ҌP9����-��
�ߠ�&=�����vl��SA ��Qf�4��R ����;��r�V����7�Q��j=�a�'M��8j07�9V�a��ģv6�&�����i�i�~K=e
O���>JW��U�PG���G�8~iw���%~��0ZUMi�Dlh�SMW&�0����~�Օ�V�� �K��������TAY8�!�AӦ�[Qh�h�4H0.j�n��j���n��Xy?f�~��h�dv�fj�x���" U��
�Ў`!KB�������طw��P#Qg+m\in7B1�h�5�@�M	E�"HA��o��i!�N���D
�7���bze���CX4���ݚڌ�[�!>��0�$y��&b0��>�"
���N|�+_���Q�#�b��7O6�ؘv����PH}�d�t�DUf"K��%�{��12<f��BN�I<��ø��wb��]���o6��8�N�<p�5�&��0�x�Ԇ�N��Gkrm#�/|�KI�p������*���濻������Mۼ+���~�����7�z3"Ѵ���͹��J���풝�}�V���y������'�zP��H@%����=�9*:������8s�"��\��v���/��ŷ���_�E�C��=-�bO<� ����O&��[^M��1xo۹�w�Ɉ���=ط{^���o]vd�b��G@]0����e!�G��Љ�����DxMm���7��͓�i��7�ar�(6��brb�c�T�i�`��><؏Q��4���OŐJD� M��D#�:ڞ1F*A��N2A4L�9��AAD%�K ��棶��Q˕r�	Q����#���;q"Hb|�T2�djz�4���0���EA�z���H�@��}:��18���{y�}�S�|��ÄEt3��~LNM�G��x������%*����γ��.�٦�!9H%�o^�~��!MJA��$�?wej�5��s��XE���A- �5�cj��ޑ>+���,:����JQ�|����A���q�~�mq���D�jRT��k�h�_���r�e,m4H�-�J�U����
����B����w��e+�Vm����Ut{P��q�D�V���n���)�UK��qI���P�v��ce5�a]H���($(qF�l@��)g��l��t^r�~��u��U/%؏k�:`��G[y����4�{כ��^��{���O&&���L� �?��+&&�n�������V]�d�!�Dp`#�S�I�q`�.j���kj�Ɖ\��WȼK� Z��>^��J�P���IB�D����a�B� �B������!����7� KLX�������v
�#��p�BJ[�Uc����%��>"�[�G���� t�/�mN�u-���h���:fϝ��_̕hI�e27;K���h �\�f��q��aB��`��US�h�F��K�!�X�����c~B�n݅���~�1�:s޾I�P~�Bc~a�ꪅ��Ve���T�d��ƿ�W�oz�0������}>����쑣��N��r�~��o����?� 1�X*��=�c����<���el�2�����J{�J�>}�fIܻ��3.2�KgNc��S�8�}��:��<l)�k�<}�I�}�����#N���F��F�( ��v�.�g��?˥f��Q���=��g�iԳ�W�C�l)n��D�t�u�v!�{e뾡S�����Ȭ�u�wX���1�F��s���N<Kˢ���^/��7���^r�v���T^K޹�]���
��,ӧR䣴LP�����Լ�n"y�#��6<<��w¥-��S�5A��N�G����Q��)&�65��ʊ��|����=�1��Uz�:L�W����D��.�S�Zx�Of�Yz
,�@��r�#ڑ<:CuRҢ�5����⬸M�n��H�̇n�l�oe����՘���F�ʫ���&0�W �0���K�Zz�@z�T�:?��k���rR�ɤi��h�����D����-[�##�n�\}�>����PC��[1�� �G�Z:��@�ݳ�~˭x��o1+e��0v�ތ��~�y��^g�稜w�سoƧ6SKIc�/��,k��^
�D"I�6�={�ar�fʢ:�ҴS@a#�2Z����`kʸ��{�܉<�ꢰ�B%�t�	 6R4F?�H�k��|!��e��˴48�8�:��|�࿠c�B����y�/����(DVȜ3��������R�P x�g�r�2��F8(�
4{ggfQ&���k���lTQ�i���Kx�ۭik]�SNV.�j�+ej�4�^��>�1m�C�:��\��Ha%Ģũ�(ϟ>����k:`�gN�̉�(̭�5�݆o�	�(0�F���UZ�Z�\\X���2�����F�ڶ���;�S�߹w&��eIhSay��o��Ȉ0�`�#�f旰HKzfu�}��9l���ؠ�ѪmQa�%��X��3���?|���?����w��_�f/��)��V���9�Z@z'�M�rb����݊���x�k��J�0=������"pe*W:�D���q����*�u*a��/{��Q�����y�}�z�6�#e@�]�n,f:(j���l/-���LE�{�"�:Ѣ	R�'"��;
�-7������Tb�|��_ݓ�k�������6F=+Rx5�T]��JK�5��ݯի`�����ޤ��Q��H[T@;�6��,��LJ�0Z2:BB�of�Fy�f|	��Ơ�	�?�~%ѳr�v��d�f�uۼJU7�d��7T��#����*p��4�ەN�Ǵ�nb��}RB�𥆆[��2>)��l��"f�,c�����k>�ML`��a��I
���D͑�c�v<���~�S��o��H�(T���h��\)B�(vP���W�������]XS�(�'�k�*N+)Oc/�K�=@A�QZB�E�>w	'N�º��X_�{5W����Db}��Bh�I 9�Wc���!� ʲD�0��ɠG��OxA"�	g2`���	;�^ر9�s�4�^�ߪ��PD��N��7V7l6����yc�^S,[5��،k�)�ju[�����������;18<�\�`�X2yY��L���%b��Ŵu�����V�m�C��T���پ�o���EZ���IuR{BiC��\����w��_�����o����]��;�'��o���c�.2M?�b����?F�?E������(i̅>�E,��B�2�m�g��#H���c��]R������l�<�-�Ǐ��_�6�����s����O[7Sçc��O��R �~Tj!<sz���-�M_0�A�A�˿��L�t��1����{���J���:xK�Y����.^��)�����y��nA��������u���2;�w���8��E�$���jyjIf��:��ߥU+\�ۘ1�M����!�HX�<(߫�K��X.��g<�4k'�o�J��94�8'�O�	��P�8�� +*(��I�ٜ����b�B2��=�zd�֔/��a�-ޫ�PXF��b�m
��&��T���[:�]�0G��Ti���k�E�VW�d�`��#A~!0��a��?�����ų4�W�������A���ӈ�4\Q/H�m.�K��W���G�̗ ec���O#�L A��� �%� ]L���T�}��$�d�Z��B�陼@>ZBø��nl�����o�^���X������D8î�	\K�59>j�ȭ���Y0�V��4	�YZE��q���%�P֜���Y7#�^��Z/�y���fziq1�ZE�e�-NA���:�<j+����g�B���v��Ue���7��:��J&Gƭ�auZ��7�}5x���\�՘l�����狹x8�����Ė1�� ��Y2r?wO����3h��B:�0{�<��ʗp��3d�u3�@�[��30>~E~��&�P-~l5h!��p�V���|��{�?��������g��_>�(�l�&A�'�I��EB����0�:.�T�M�'�٤GJ�R��JlD�6ֽ6�,��qt:���8�z���Ob��02��y�q��3�hh�\�)d�Y�g�H���T���w�'>�~L���,,ۮ����O�cؗ�?'Ε/����^|�?���2�\/g�����:N)����s/����^�Ų���{6���i�����;5h�l����ژ�o`��>�#*�l[�R��Ԏ'��e2�Z=�C1aP�L�.�	��(k�ID�)�F�tV/����xo̼��������Uu�j�&Y?��|O��M�& ��6�cG��i�X��K��"v6i�+�آ
	HK�)�#�;�=�Y����ńF�H&�a��Tw	�ȫ{�R
�MImb@R��jBE@�QS��?~Pe��E�=��-��B��B1������r��l�� �j���F���JfU���C�<5�8L�;�Q���lѾ$�ЇJ�L��A���O`��'�,����ţ�S�Q���"6�"a��l�L��-W�c#����ryZ$,��U4.Q�xSb9��i�<EN��:�U�KE
�&-
�by����j|�Q�-���"CQX�øI
�͛'��E.����X�\k�ʼ��IZ~�T��_+�(xZ�the����C��[�՗�b.@%@���8sr��<l{뎝��x��{p��'p��1<���ҟ�W�z같�2�g��C�cxxW]}���S�u���� �Y�&�iIrY
�"r�8�}���}^��w�=�0�ſ�M|��ny��\�c�B-���Zj�
[���i=�A*��YY�h�;��P.��NL�޲�;�pmi�Μ���3���%;�82k,�z��i�1�����w�?�A���u��=�a�wa���<�4*��3��,��ΩJDؾ}�ܸ���0L�6ڲ�����gm��%�`�����46yp�M{�e�~�����i	S脣�� ���j�:�m���Q =�h5Tdw�H�R���,I�lw	+�i(f��}㋼ZQ�Ҙ�ð5u��sϨؙ��P
i֘&#0O'�һ|��i;?�i�S�W��Մ�s��O�����c]�*,���z+٩�F�v�u��c[c'9�{K�"�Wy��pJTy�Ǌ,'�vM4p���2��0�Sj�	P�r�%�1�%�(����T#��ή��?�l#�;q���J����%@��Fbp��gi!iӉ��q��1���Q�V�__'s�Q0�O4`ݑ��W�@[Ϭ���!J-Efi�������F(��{?�Qj��i��J����r�L��;T^�LT+�(ՕWk^������XWYy|�R[���[d�
�,�u�Z�ul�(�PҞ--�d�����c>*������r�#�I�Q����̫�1,Za�&�'�-�#	?�ƴ�'�H���%)��N���m�}=±���/����111���{h �����7�{��-4�>��uo����Q�`���_������Wￊ
)԰��MN�SyP��W�O?�8.�?��g�"Ea�s?�^|�;�[������;>���韥E����U�y�(��1s�,N�9˪�X3j6���"�:q
ǟ9�ť\8w�N?M�Y�S��}܋c'�Y=�WVq���n��J�
Q�kf����w���_���߆���xխ���ҩS��l:�}73��/��q��������K8�2�k;�Û�����O0�����S�&d�4FG\�4�3�y�
���"O����]K�!h߻2y���b�E30'F��pc)��zԋ2�ێ���>"	��i�W]vΌ6���(�b��q]�)^� �R�+��/��gu�K��n�MF��`��n��$���|/.f-'_'��3�ٳ�ȉg��HS��=��'��Ŝr��+˪�R�yK_|���WVN#aV 
y�G���g���wN���

��࠭`0rYڳ�N�>e6i���F��TQ���[����Q�ס��$D�P3y/�T�X��%˒x��r�,�c-3G�1�?��-;$����5��k�����s�X�USm00:����0b��OA���˳��@�dڊ&Kt��+�D8M���Ѻl�M�q�G3	��}n�ߔ���ۅ{:��G���ڰ���m��$�����H��@�m��1�|!�|�j,G�~KKKN����;Y@���$�։�
BY;u6������{����v;^K�D�齀#R(�Ӵ:K�G�~��`j��m�v�B<=@�݋ki�lۻ��_������S��{�=�����bӖ-�!��yZ��ė�@!uaڎ�x�'p��)준{�>�M�S�s����aV�����XY[���2k�8�Н8}i��_M��ª6�j����i�i�d���G��}�=�
�ES���<m�1]{�uFc��5�%�y�vZ<���7�D:��{~�=عg�Y֚E)X;�\�r^v�-�،�g�q��c8Gkj��8��{����m��[(�^y�-�'�����i�����Nݮn�tע`y��w�O|�)��$��MSG�
��0�4��v�_Yӑ
%Ե;=y�bg�:21�4Y�1�a�V��֔?�X�D�@I�j�����Nx��Abnhl�z[���~�C�My���M@8�46(!gi(-�����q��bL}��9��z��QW������V�rRp�;�9\�	%���O��c�8�z����c���;��ɘW�Y�5)�:�G?��;�,d�o�@�ؠ�	��Ye!B^2?Α���4/>�,5>]����A�!�D����j�D�:��<p��B�?��T;Ƈ1���^��U_#�ͣ\kP�R��O��Z��8�ٷ��R���c(e簰�J�5�dz����&���u�ҩ>ۭxyq�v���,����"�EhjS�e���p֥H/9���d{�t��ӹ<4��U$XƗ�Ɓ��3ᘙ]��֘/�)�]$y'kS+拥
��>��r�����tx��h�MS�:�ٮ�'���W�g��^�ؽ��
x��s)~���B�ͩ��=a늆��ɨ��oA�� _�=���p��?|;���~�_a���L:È��e�$Buc<�$��<����1k�7�o��'ÎR�{:X�`�旿N%%��g�c��94qۻ~���ċ������nz����|�V�1
�,�	7���֥"�moĻ~�')LwҺ.!�b˶mX�fmA�5�]�WS�j���,	,��LLN�5��o�<L�
���cGiU=���u����7�oy�[0<1f�Fdt���j���5�[���n#�]�#w�9�SH�:]O�1��?���1*4q�j5ll䱲Z@��B�Y�B{�~
���7
�;���0���Y���v'�j��Qӏ�+����vE��1����=�	K��(Q8��}�;˞M ���/��w����}�Q��P1[F/�>!����i�¸)PeI�܀���	�%��to=^�tzw&|����b���鵧�1}Y��t�g�֜���}���#>�$|�u��#�D)|hvv�t�d�ڰ�E��B�եD	
M�N����ppx Wm�ö�4XՍCL�Zd��6����I ��k���o܍5��Kg�MlP�eCR��W|����h�1�j}!l�b}�fΜ@C���h�C�݇hz�7O��][112l���qy��kzf�C�B�mJ#��b������B������R8Ԇ��F�mS^������1�kcWj'�܊�C�H�RX��[Xfd����=ש����o�Ē��q��Y~QCұ]��T�p*�R_��D5���ضu~�����LO�|AG�Ri�g*����&�����'p��Cx���#8��C���w��o|���WQ+���ݎ����p��7��tƖ����Cz��q�X�:=rb�&���������x'�<���ͤ�fj+	����aj�5��Moŏ��{����nڎ�Pؽ��o���Waj��Tvv^��_�F��{ރW��5�Ŵod�n���{��f
���e���}��֭��R
��q*&�5}֍p$��MS8�4�m�D�>lٲ	;����o�z /��v��]�d�������8{p��������!x�ѯ����])�m�O{�S��~h������62Z����g�Rˣ�o�
j�Y���2Z5�V�v8��+���v uZ=U�PqG�p��Wм!�pܡcY.��r+�.E^Aﴔ���4�aE�L�,c������N(��V�LZX��)>���SYD�~Қ&��C��pJ�Q��DU��<�e��^�P��f}�U��i�)�xUU<�f��^�0�%�|��u4���]w�|�>�o?�l�V@�1B2����j�O�A�G��>�E'_�;H�GS����q��k��Xڃ�ɴ
k�m�(�
8����W�Tn�[��c?�*���W3�<���/"?�@G�/��2�`���	����3�E~���P��q��I<u2���v]�R����q��;�u4���5���ԓ��;?��	�!t|c4~��<���0d�5"�fa�[�A�u�������(|�y�&��-H��������O�Z����]xEj7�؅��'ʵq��e�b��mp��a]�=��L%�5�P����¿����Cާ�ְ��BF>���N-��a�/����������B��Ez��)����ef�:��NM��'���q��Y��
s��7>��b�����[��N
�>⑦Xj��.,��Jv��DT(�0���z�b{�C!��⃻F�����7-���pe�i�q�d:��6�$�:��7�g�ʪ�vR�l�U�R��ҊSy��I	�U)Xڰ6��ƈx��Yߙ�`lڲ��4��P�ѓu'0�jC��Q�R�|�#L��2Ktj�aS�	�������v:R�Id�?w�/ߋN����Z��c�q6�7nV��B������)����]��{�}O<u�@�/Z~��
D�F���j	���6���f�z�v
��C���{g��,	1�ciW��5��
��h�6m�kzu�۲2o�θ�U��巤(@�c��J�� <6n���V�,]�%�V�u5��rm7�Z�H�B{��IK*��^���Uv�Dp�כ��0&|Lѓv��Z�<�ͺ��kk������<	�E'��z����㎳|��S�j�,D�Eg膩�`5�C��&$%�Ĩe��eµ�g8�����8~���-U+X\�a.��rуT4�[l��@3�8q����/�Aͮ���a1C�Q�ВI`<���.�.،��*M����0��L�4���������Iu�,�f�3�:Q�������B�8�e�f��L�mLM� ez�u'ڸ�a�X�'����T\Ǔk�h���3�°ۇ��a��&	� �etD�@�(��!��=!���z�ƃ��>����Ο��O�=�*��3�9Sh̹(c���~�����C����d��~�o
`a4�S}�aZ������/}	^�ڛ񆷽o|󏘦�c�vĢa��.8�c�+2��YgM{OSpk�N?���N]%�*"d�t��A?5�h	�y�
�,3�PM��8���ʢ��ꦛ����gfaZ�g��Yv=+��sg?�p��8�gYe����Q���Ŝ����._��~��W�.��ئ$t��	����7>�?p���M��[����&s���:82��&��:�/�/bzz�K�(e�'���8>:��X�v^&�+�_-��)�٪�ۏ����+��
��;!�Ѿ�;v�zuxiF��dq�DSsHK��v_&�Ĥ���1��]UV{�i҂�H�=���N6�H'U��������zgr��jZ�&?8kx.u��{:H|a9Xݜ��Q(�i��Ƀm���z8;��.�'��Dax�E�X����w����W>��4�0�"0�m��i��$W$2l���v&����o�pri'�2X��p)W��K+81W�@	P{��V��JO�_��Km\X���\�85˼;>����g�U�,�u?ίp�|�uʈ����l�B/[Ʊ�*�e�[�#�\B���R����<B		���Z9K��Y&��|�/����Þ�4vN�i�X*�㱥c(�ˈҬ����wB۶lf�hz�Vѩ�|B̏BHӀŘru�9v��TÉ1j�G��a���&�R}}6�Z�Y�+\*��M/�ɺ�~�'�{ݭ�x����ðA���N_���ȝ(��"�`P�Oaׁ�زc+���Q�n�^�O����!�������s�9���;�8�p����ݳ���x�w�=�����k]-��Q�����=�����^7�y�������ޓ�9�}~��Q��G?�0����&�ٯB��8F�8��%}Tr�d�nd�3��y�Vk��"d�	�Z����z� W1O]ʪ��"��טO�-���*�N����[х�-z�-<�Pujɉ)I,�)L]:�M}dut�r��8����h���Gs���Q8���L��ԑ��md�v���wb��{3q�睮C��th�W�w���A�g۳9���z-�I����
�3>�F�I��&Ҿfn�Ť;MT��W����M�GN���� K�3]*�d����3�&.��1w!�Ŝ���ܬj X��qr���*�)T���t��*ZE�Yg�BЅ%�~���:"���X�Q��VB�FË:+�x������,�)S�6�4�|�������~b!
W
�\�d�h�N>��c��l���)lI��ma!���7Ρ�Y����O��m;����(.�^�ڱ���D���[k,����̷l\5��1�㪃Wc������Ν��g�>Z9/ǭ�ގ���x׏�^���`��ݶ^�%Agq���u��L���g�N�?X�?t?tߏ���f\$=u���k������� m��6���j2~�6J�S���:�@8@�������V���b�Z �(�D�Hzx��E�a�vA]v��@�W��i9c>u*��dL2�^�w����������������z��{��EV��R�kL�t��^i:]� L�1�^�Qp'>����/��`J��;E��?��R�kH�q����.L��@�ޠUȼ��m֙<Ê?�\n��5q�ͺK�I�w
�&V`��*��(6�?������\a[��x�**�*�3%,���<X�j/rE
0�vH�7�J��Vi�t@��R�*�+�a��Fo{;��
Y��(w�l �W��Mz[��c����ׅ�6�ԞF�(:�$:�����Q�j�]�rBX\�J�����7���Z���yt�	#5�%�Jٺ(��B��1r���jf�?���L�Cm�A5����q��yoW�`Ї��Q\�5��w��ׯ�2~�7~����o��W>��z�O�/����(��Yʣ{�9KCBQi:�=d�����?�Ć�4N�m�r��(��bm�,6�tG�!D�4K�#K�^���N�V!�w#����v����f��:����XZ_���
ʴv>�Lʠؼ�9B��F(W2�.=�~d���Q\�z�k�^��W��W��:�{m,~+!B:'��P��h�ǧ��'q�8�/�[!_��Fi:]k*�x�<sPy)Ȋ׋s�t�]�u=��Hҝ���Q �n1f�9u3ަ�[ 	��s7/	!B��Aa�Lri���"(5�d�u+��4y�5���,�X�dx�qg�kc)&ᵚ���\.?+�3- Ĭ.�3�Rzӊ��2A< W*wF$��G����3�+�]��<QZi�!�"��1D^�b)�baSq���\����@�B�QT�^��Tf>�A!�1�ӈh7i�oeЩN#W_D�U��q���zyZ~�bK3p�Q%1�xr��V0���sN�:��tk	\.�!��b���ػo�]���c]u���;�u�N�=a��9�L�������'N�\G�)���C%�^���{00�F:�i�>
��u+k�X(� ��G+�d�d�&�l�S��Sj��X�c�R�;�F�o�f��q�����#�S��h�K3,�؈B\f�]�����.�F����?x�𬟂k�ܙs|��"p�v_ЦS^)�MB�i���5�od>.-�P.��u�p!ouƳ���>� �����%��F�4we�g�>׉Ո���ޞw�,g��e�,��#�=d�::@�NY)������$w����(��� �xѠ�Ck8C:�@?}�G�>2wBH� ������ <�it�Q
"j�t4�;B�/צ!�&�`G�v&I:F�j*+�7�Gs��a`���C�oBhk?��)��!�sS�Q�pGiV��Џ�=��;��G����d��m�e�6�m&�a0fRQ�A�u��,� ��V[m��0�"��ʫ"�k���,��[�9�sOއNvV	;��ȳ{�9���p�����MѴO���F~�a��z��99?��W��C�C�9
�f�:r�`]���K���ɏb��=�0��_�cH�6��㳞�Z��t�L~�ծ��ؒL��{�(�^��t�{(e���L[:v�8��e��\I#�Q��n�5�k��h�<��Q���ime��G�Ξ���JqSe4�wDw�W���a��hy�8�v[���0�L7�H|����Օ�]��Y��s��t�Y>z�c�Ǯ�H�����4�Ƽ���$]�s��U��D`�(�<�ڠ�����:��G$A��Fm�"��BI"��1W�a��iF���)�N!42�ؐf�� �7�X,��T��H�B�ix�i��!�y��aD����QsE�n�LTl<lO��mG��@b�$��鋠\s�j�_)S)DF�`ޞ��a
�~4�a4�DV��2J� �O�Ѹ�oAIc]����0P�jp�&%0����0�ߍ/��y�P��t
��<�V�<����N�N�נrW��	Q�|g�u�����q`�t-�g�S>����������	5�8(uX�W[��'%��l�W$��LVO�B�#O��!�m����X.���F.!��ޓ�}�{� ���E�����WK�����3��pؙ�$��<�<��6��a{�q�[�Io�p�Vm ܪ�oV�ik�f�IҲR�	�L[���?m�[�ב)�m@O�8W	�f�G9���|+o�Z��Y
����Z��Y&�S����^ν�;GB�W~�(?*����i����$�A�)$�5�/3�ԪC{iYג�Ksf�uNw�Em�a��2�`�z
�G�ܣT�-G��~mX�w�'@3��-� �I���0}�8�0%_��
U��}�h,�f�uB1���XL�������J�����7���i�5y_����u�y��sΌ�.��JL]���Ȩ��1
�`�cV#���@	Z�qZ�2�fU`g=)��SnP�u,�_�����Y�W�����k����p��t����������������7g�����z�b3�h��:�V�cdj7���h�"쳉a�	-�И��|KG�Tȸ���=-)�H>�Q�m��"�y�N�h�QA�������0��y��\@��ob�!
��qm~�qȢ�w{ȧb��ӷ����'o����m1e)�������`k��"��b9��3�Tq=�CQ���z|B�%�l� ��y�1���>�9��{�['I�|el{iι���	{���Ђ<2f�,Z/T�m�-Y�)h4�C�ռ�Pm6&��ݠ�S�gM�7�O���>�ƬIO���[���� 3fLD3$|��g��?X0
ީ���o^�G+��	l[d�:vZ[<�h������}�i��>��rR;�N��5	"�����C�l�`�*:�g�C�	"�GjQ�Ghҹ�:�S;��Xi$"�-Dl�����̏Q�q���~�.d.>M3�����g��W���5��@�?�	��w�Ӌ�b��미�p�	{����q%�� RF:K�9q��0�<�o�m��zg̣^ڜ�-yިӾw˨?�[f�g�,(��&���#�|��@���^�򳥤L-c}r�n�ƕq�u7X�3�W�.�7�pR0�z;������w{�F�����-*�oϖ�rQ׮�9u삣X�>�����&�_/@���^�v��n�^p��w�+T*yK��W�Ga��W�URρk�^��]�/�Q�0:��T����{:;k����%<���p��#���T^*�^� y��z�iG}�%�V�:HNZ:D
?�`$A��S@��Q!]����gi����L��#;"3'�Qx�h���|�%�����r���T�&�Zǻ��U�!�#V~���:����K��F�SP����5,��
����X�m,��� �rƭ�Y�)��3fml�|��B�{�^[��;�vL|�����F�{��Y곝 �{Mfp�3T{�Xxf�L���봶U��m���d��m Db��%v��#�(��&05���(t:e2[��>�����&4=,c3���)�����4����4%R�u�i�Y<4�
�6
� j#ZN~"�*k^��V�����i�P��G��Qc��Ӧl�(4t����T,:=/�n�B�@���J(W�Y�����]�m9��&��<�X�(�� ��G�ul��L�%��Ο=��O܋�SO�SYs�ؼ�i�j5����W��`k?]�{���V�+]�"rJ�a�|�O�!B�<�������t��^v��evXQG��J���w+�b�&حC�x!��7C=���cCͷ����dc�o,�e�0���Oߝt�x�]�l�N��k�E��w�?�'���)Vv�3�Ъ�:;i����+���r�d�J�91TѬ�qrw��q����`�M�>[���6���a�����6���������p�ߘ�ĉ�:U�S~y�Q���lm˯�:ӒrU�sɒ.WѪ.t+���,Π�9�J��i4+�Ъ��ϑW,��L=C�e:�QaTE�~+gǥ�W��4�މ��W8{�	D�!;G,"Sl�Q'��r�u�r�u�iU�S2=�����a��y{=,?�^E;�h
���!-�(�����p��>$i
 ���jr���P%/�R.��Ev���x��^;VW����H��*�脆P��Qպ!*�R���REr�<�m�wBO�m�����%�C�� ��<-g�m��h��.��[�s��t�Y��~t�z5�drC���m/��	'�Qs�~3�H���Zmw�q���{_��
lZ�gIT�/d�Qα�hi�O�����F�c=�~��R���6g�J�6�C!��f/�Jo@V�)�|6NLHu�jЏ�M6�vS�K�O���m��`h&�[�y�0l��*��P��_�3���$B[G�<|^7��%!��T#h1�P��M��iv���?���x�-�7񕧿�O��k���>��7�����1���F�>���3�l��ؓ�]�����O�,�2a�J�cl�&Ć�"��G<=L��F7�(��R�)M}ы�9m���{6���]D�?�w���X��.��1�Ep.�O���!��7��6e^��iL��QD��bX�{	�����A�l���Ճ��u�=)k����pB[���z��EGyCvf	���1H0H�KT����΄�$%�W�nJ%a;(������,S�Q#�sb Y������.�J�S�BFM[
q�nL����I���U	�L7��?�Z]�D�[�*eS���w��V$L[{ȉt��V��=~>K����	 �*ҕ�:-|u���m��`T�t"�pQ㻦Poj�`�1��z��,���mS�%xT���YO��V��Z,�I%�A����=*�6 ��YFƓ�e~�
���
i�uD	��0� �[��&�h{+�F�P�Y[�Y�K��o�^t�H�qs��l.*yK���3����(�?5�C�j�W�*��g�'��%e�ȥ<�Ƨ��K1��Ϝ�c>�GOM�ha	�U�bA��������a�VO����?���X�$��g���]�)�.�ob6�e��#��ƍ��^���jd��h�J��,�&k����656��g[SN�P�_g�)I�����W���0"9~u��) �y�O�wK̶��<���O9GA�*u�&wx�f�5�y� @��6�4&�ˤ� ��p��襋�ʼ����i���v�Σ�x�G?��E6�P�tCi�Vq)�B̈́"�O�)�Hx���e��"rim�8�ͥ�;Y3ړ��Cjk��Ij�t0���'�3n�Ġ�,TrVX'3Ҙ�lc
!���� �46�?��^{��H(^�C݀
 �՘P���b�^�����	Q��X&���[_u<��v�n|z�OPieX�~|x���W�(�w���%M��6mGE<���hT�&�6q�
E��/Q� Hx�´�)2�$F'����n;�f��hم�>jT��.�#�Jb�ǲ꠹��&���	�PHUւ
���a4�K�"��g�k`�)�İ�n+!��������$�H��C�Z̻^k�ʺ5k�""�����ե!+zR��Gi "6֧E�6�	H#$U2�(f��HQ_��&A�hmf�f-��,,�3�aB���mH�B0�VN�C�Dc��X�2�#����Dx�_���$VŠ��$�Օ*� :�Ȑ��a�Z,_8�����4��a�{���	^j�:�X,��H&6QG��g7���j� �Ԭ;d�6EVa��d��{��h�V.!���#�!��jd�!�,*}~�ǖ����F6������5��5��\Z�ˋT"s��:JH�I�J�0�ݟ�\�#F�v�2pQ˧v�|���)�	�*�3Z��r+��oh��Ґ
���W6�`@<g�<L/��G�
V��$����`�^��뀔N����Eǁ���
���xH3�"��D��y�!��}���tBm���mX[C���^%�}��3��8iIB��Vw\����"�$�t�"�>�g.��\a\h���&1HMS�h�ov���X[-c�8�e
��/N���ݵ� �Hn���C9W2�4L���	����N1�&�D$]>*Z�i�������o�Ӗ���VIg+��kPY:V�(@¥�KW��vUAD�/��g0'�SD)���-i�)����^�����V%\��@G�4yW#\Z~
�-
����簲D����A0�B��r�p|�P�BD$C�o��������G�K�ҒV%�H�R�W�/i��� ��V��xdAxC5Oګ����5@ICf��3�("u�G���������#����(<��Ƭ'�C���r�˧:y*|j��/��*.+EnA��>��߲��%$��������GTPBh
���f��o���ײ!��o�,6�T�<y�N�dbd�@QZA�a��W���(�$���H�R�"G�AXHS�ux���B�'F��x.;QS�.jx�ӄ�	kfGg��&�� bzb8h�b���(T����M�����G��m$����v�f���#\�B,i�L�J�Z��)AX'�4M��[�t鼢X"im�T�=ˡ�|!Mu�PxQu��Z�2�3d$-Z��Yoխ�2����:�X'��RmS@�Ơ����,��H{��"��\��K͊yK����l_?��V2�O�984�d:�*����*�Ō�"���ı�Z�8*�!x�خ�˳dX��"K'0��F��Q�h��"	>A.3�R����֧f������,/�aya�f~��ȃt\8���7RPO�V^�e�O ���Pj"Ca��1��� q�B�QE�į6J�&l��L��yN!S�WQ��ba:�S�Q���� �L3V5����`�j��&���a�L�Y�)����P����T��d���d>�� -���´����T�%l���hZ]a%�t���;��m�6(�#�$�����7M`��	�0�9@�YE��Z,��%r��e��H?i�Lu,=���v��Ґdr����-,.�̹������K�k/b�t��a�S�z��,�k��.c5����6d=CRT��$Lȋ�1>�CM�CR�H��faӦ)�������%��=�ݑ�-�ME)�cn4�פ��G�H\'�HWw���-�du����kݢ�H�eb*����_�	F߿��[��ˊ-�)��f�������Q �ɗhxhM$��+��|T��$.�6-�F�����x�/}��,�f2�4_܃A�թ�K!S�Q0��[� �����M
�
�fƄ		2jr,��R�1��@S��$;�i�,����%s���@�d��ce�Ek���Q�*��<*R������n6��-��Mbt����5���8<�Nt m�����N��*d�f��A�L|����7��P����_��;�|-���~g�Z�q�F\w�VSau��ja6x>S���"�dI�K�H˶��ږ%$����^ʸ�AZG�"V�6�򪭨��Z% 4���ع� �F؈�/��
�`.��]���"<�d(�4p��!��}����B,CN����Fk�BF�n�H4L�PC��Fǣk-��Z]<: P���%�d�2�Ӄ}ƤJ�|؄W Ėb�Ą�mj�����*u�b9"���A�I�Jnu��Iu!�&�B���LLBE�8�4>���P�%|$E���0��)�>����du$����FL8���!Km��1w���D�G�?�vr�d�m�F%����O�3sC��M��,_,Eش�X=���G�?S�5\����?���d׳��e2O�+�*�S����%u���X*j�O��K�҉>��Y7��NZ5%d�{���Ԏ��,"������fSF�,�Z-GAA��%ɛ6��2^�$z�Z��R��%�mM�mR/Q騔LaiR�+h[.
��v���P��$Ec�Rƥ�I��S#~�D�l�$��,���v>ljL?pہ�)-<���hm���9��үݢFk�^��KAH�W�p����(H��Ɯ���5V��S ��p��%�Z��\}��:����b!*l����e��	3�)���`&t�*N����L_ʏ�c���<�7TXqp�_TX��;�_���΄���1G���4��&��/+M��J "�7|0��W�:��X^%DtoB�i|7�WYGEc]��DoZTZ$|$c%�l�7�:5Re��L���u֕ʊ�J��'/����i6M��'2�<%!���ʝ\�V�߄)��W�5�Y+3���aJ�bc{�W0�"�7ͼ�,�Ԥ�J�w��U"��G��駕5���j�,M���-F�'��(�|�a�H�u2#�Z��$Ou͕c�m\d>U��v��r�}h�ꛗ�"�D�t��0T&-b^����>נ��w��wq���P��ќ�S��`���n��.�Bj`���b�q$��X���r�k f�Y�� �P�IhHk�0�X.i��2�Ҵ��4cG]�Nw�`� `��F6�����O�#S�b:#2��]��O
�$|�n���D�B[ic6c��K$�hdH$:%T]�����Q�H;p�a��b��l�pD]�n;%R�X$#3��e)<i!u��K�q�L���#KS��Z�W���V($`�"dj(v����\��Dh�&l�;H@�X?/��VMr�Qn%*"(1�D:�t܈[acy���̳��C=<L|��o�[Ϣ4�������"�O�"�s/�~�	lm�T�@��A'#�r�nH�ϗut�UV����:�D�6�����EB_�}d���n�ZT[KkG�o!����|�l�X��^;���"Tu<��h�ĽJ�鎶�#��T\^��n2ii��UX)s�	G���ḯ���'���nQ�wu���y%��� ,��5GQNXk�LL�Eda���Bnu3���M^�It���%���@�����a���ב7�K�a��䦞v2��+a��R�<��L�P��C�45Q�J-�B)K�M>A��V���71�����:V=X���f[��J�cz�b��:��nL���%c�"�A�cou�������UK�8�c�Y�!F�zW�0���U��Zo��D��͐R����L�h�md�E�Z��0���[��"'�Sߜ�	�>|o��Ǚ�I-)#Rh�$Q�� ��!5����u�0�S����)V[��?y���"W"����HT��Sd�V�,��"�B�G&�ce��ԦvZ�t�V�1
�5�	�v���-�֨��4��r�@bH>"�6���b!�>{���]#0J+��=A�q����o?�C���$�[�2-���KKu3�A���I}Z�U[Fm�!tV�B�Q"#Wc/A��O�t�J���,��U&�����`��<�~�����7�c~u��?��~52Mu��=�v:��� �	Ӣ4;jj�ߖ�nx��G�,@+(g��Ǻژ>�n���2�����Y}g�p5f��D��Ƶ!Ҹ��h/䬅i³Q5�!B���B�Gت11W���t��?d��4��N^�!a�b�Ŵ�M�F��D���L�1�v��!{�~.kVk�Zd��J��|Od�!�R*�xOeP��R��I�)\���uj�p�.$��AZ?�� +Ҝo�*�}HP yb>~��#�P��X�#�#2!�F֖���q�XFY�Uj��� MW�@�7H�22,�V+7P����UP���	"
_D�>!᭠�>������c\d�]��`]��y�YV�[��>T����MF���*�y�&Y�X��K!�85��U�2�v)
��.���7u���4��OXI��O�HK�q��G����.T8����d���h$�=���!���8J|� r�=�j5�TWx�%f�4��E�X�m�W���K�i-e.<@jQ��xA!�	�r�����c�I3��`ôX��Z�QY����=�2�(?���/�%�JM�H��<I�Q)v�V�������к����b����"�/N��O���%D|Ml`|d��+�{����O�W�H3�>��QaʕQ�F1���j+M�#�T^�G�O�,�6���񉷨��C�JS�%`��f���e�j6 �ԽzvX	���꨾Sv:uZ�A
n�h�6�JK-�l��A�П�Ԏʴ��Ξ����L�х}�
���u�O�.v��Ѹ���s��
s���F0xX�$	�_�M���5x~����Bw�ue"(R��h �^l�ƚ �(d��0��b�DA�C�����i�[+�@!��6Odu�STChR�d�Ǫ��Gs�t��j$����B�Diy���T���V� �C�M��5���$��20q�A����dd��-��i��[��&&f!�^�K� X[i6Fԅ������@����j��G��:R$�0
ddK�<�u2�6J���I���u��I�#����s�q���[d��b����/jv�]��cӭiq6�ŵ(�VJ����3M���C&&��.-+�ӖD��	�@��d�~��f�Rf�G;@Dc����4���A2MAe\�� a��i]:��N0L�B'B�F(�t�kJ��5�cڔ�'J�#�-��KM�Ԡi��L%�H2�8	����0Ђe4����0�R��~j�j��0��T�b��(�:�(�d:�(���}�����'�4KH
K�p���6P�h���0����8���S�lq_�@�6�[5�(-���4R�u��m�;5��BmU�}�<���,Li�^2dM0fD�ũ�G��:����p��|�u�a^��n�H<Űl?�4a"�A:FMP�C���8q�J/˴��:_�R��f��Ug�+�GL�v/Q��x���d��!�A���mL�	?a�=.X�-Ĝ4sOʆ��g�I�1ID/�.�>�ѫ��&(�}���w�{Y<*G�~u*rH=l���
���1lٹ�t�Gvq޺�%̕��3��X�W0sq�>�'�A6_D��B����h�G��Y&9��e���i��^J��h��E�Z���5ɀ�������ޘ7��^�E��]l�F�m������n6	��Ϧ`�a�*���s�1A!��7~҈�M&2��м�p���p�����z�3A�MҊ��Wl'��m��p�YE���������-*�������*� *S7?���0���|�w�qn1��}�$�DVW��K�FdR7�r1�U��-͠a[X�ԈZ�nj��E6Ad޾]h�cDvVH�@O|`�!iU��%n[e4v#�#�	�M�%D�9$Ҳ���
��1F�VE��j�J���� ��t�М�$aǆ�D�B��Jk��-^3�`hȴ �#,���v�讝��m�$��:zf��@��	4�r4��5�^vЋ��|n޹3G(��� 2yZ>Z7�ܪd�R��^ȫ��N��E�T#!�j'��ukk6!�Q����m�!��1��E�)Q�S�j��>�4�p!��y;f�f`թy6H\�Qe��d
����#��j���т9	�Z�B�x��Za#r��,
�\}��uZV��I|h�Yh+���Ҙ��}S�����{����7��U*
�z����e[�hd	�ȘC��\�&U
	����kJL҈G0r����K��Y
>6I��(Al�����	o4�TX��n�AAw�N�JW�̖�O�l��Q�H����#�V����q��HP֢�^�)�!a,�����j�Ci�b�^��	wՍe��`ر�¬�qD[�4XG��P ��"��R�Q������zTu��ٞ�&��F��ք�'�Q��zj
~�ð��5�CR��ۑ��.�
�pY9��1Y0vx�h��l=��f��譭XY�~
�&�/m�-�P��*��t���Z�u[*V��n�f��d�,΢�1I�!�J֓&�ԛ�Vs����'q����1Y-��6F}-�SL����rc]V�Kk
��e���g��]!�nk�5��7v�������3�cL��	���Y�턑��c^�����F^��=�2����5QW׏^��,�P?ű�5}캞p�8�%{'�I���G��������x���6�S%�N<��o�*t�%z�ƾ�e����>v����r�qT�xZ>Z�+��H�y��4Z��jAXZ�OkQԘ��Z;���I����0V�na�Rz�=K�1US��x+�n'M��F�@'<iS\[�^�8`��X%�B�a|;*����*\�<�!��O�oiZ��y���iT$ie��$ o��|��2�kv���yq��{0]9�$�	Ӫ�Sk��P�DM��έ����_�-�����Yt|#H&���eԮ�Xj�,�������&��N�>�g�Iұ
Am�JbVٜ�)bb(d2궣�P�֑+�+Mp�"k "��$Ӑ�lM� ��1����{�,��iZ��Eb�z�$�i���4��ִ�u�)�:�Yח�n���Arj���f�i�
$n
#u�LJLG*5�����,����L�rE2�B��|�i�~	���o>:<L��
�2�ט��X4a�XO�X/	p	Y�j�*uƯ�Ze�((ɴT?u%h^���sQp6��Ւ�/��n��G(�YY�k�����o�iW	Y%�&���0U>"D��`�IU�M�Ph~њb�nW��T�d,����p���{�
�M2eqP8���;�0���X�)��E���+�vxS�;�bJ�I�hw ZV%�wʶ	�i@4��0�4R�g	WmC�:$���je)��{*^��M��Wٴ_Zf�l����dLi�*E��1<�8j�R����%d�Vl\5ϫ�BE]��2�S��E�3�k��·m�E1�0�#l�	*I�*�)�fu�$����2@�	�r�4��z5Lz!#�70�\�������L��r$w�7���#ϰ
�q!MD1�wt�0Q�S�bw�c[I�Xi�Wg��>J)��s�*M+]O8��BOr�;�`�Z����/,�#�,�d�(��ڜt�#��oM�)�Ed�z<�om�������r_��	����T/DM��R �tj̄����fZ	H̜�W _t �Ƞ�l$�я���Y0�
,�~H��� RI;sS�x=}l�q :	Wt-��Gf������&������<U-�� ����|DD1	"(�i��۴N�ًi�Hm�}��{��>�d�B��}�����)k!W��{ܺrȣ�xo��KlA�_�=�P�� �5�N�xGu4x�b�͂� ��C�nu=D��ʃZ����^kF�����,5UCT@��1�
��li��9T%���F�'-
s��h[y��u�)����h��zu\�l5s+�p,
_�񚚠@-����O&��u)1|P�iɼZ�N����V�4b1a��(�g�t��/k�e�V-�B��j�����k&@[d�҅2��k�|Y|��f
i��C��_려�SPؘ�Ly�ਤP��Q`��0�,�RN� ��!Μ�V�\�5���|����;���cG�ICr{4���`�lq���ZR�n(#>��e�uu(�Pט���_�yQa`�6�Є�3���	�\Z�����e�(91r	/�\��WWj������!z�Qx�z�ť�;/%�6�T}LxQ���So���o�g֘Z�����Oc��	�nmw%F�x����B�|U�K��#�/�n���zj楍]�![T�l3�jv�Lp�5�,���8�Yb��},#l�F1��ENK�婲�b[>��S��ӽhCL�F��+T�+608î=۱}8����\�#���a�M���q,I��T�᪸��{i�Ǵ��WBZ��#�;�`��U�iM��a��<
o<�����(NW�@�gz�`aa���5͛���:i(K��諸5��s��=2�s+��1S+�^�;}V�J�g��+��;�iF� ��S"�%��Zyu�g�c���=���|����b_��$-f�Auj�� �1��M�؀�:���\��f�Ћ�Y0i��R盓�4��*%MK0���^�DX~PeE��Fau����R DЦFgۮ�A�� ��T6���JWkLdE����E(8 �ŘLDe�I\�/��*��N��*D؏붤p��)�w=�e���C�KP]�f��QdYS(���0�����$���.����:��P"C��E���$Hi�ͺQ�dX�-�e^�01�z�H8j��QkP��}'��K��J]������'"�]|�g���/

���1Me-�%
d",���Y4+y�E��D�!�G9��8��F����z��4���cYuԄK���Z0���)��9�R�Š�Sx����!u/�� ���'�h��w�B��k�Jd�)ʥ�P�.Uu�Օ/�*�K[�hZ}�Qf�j|'MX]����UŲ��.��5]���1&+����z��ړ��z��+M�̫[�A�Ǻ�������PkV	lMO��YR6."+�8�p�YbB2с	����d]���Wyl�[����i)n�7�������X[{3��;�����*U��h�At�<���63R�.+��8��TV�_�uE������z�@��EAy�RXF�3y����lf����ޓ�J�Q�Q�lZ��J�X�8G���JYa���㎺JY�.u��7� �%�ܘ�z4K�ʹ�Nl2Å4ې8�=k���g|S��n���SDZNzM�A����k�4�Tb��,��%�|�K���6(x2.��h2iu>����ʋ��w��A����(�	6��D^����,E�y)����*�*8W>�=�?o�t��u��zE�%��t�˩�����VG΄[/���J��]�B�to�%�����"3D6ذ�&x����W�(Ɨ$A���8�����/b�Ԁ+�G'����Щ���6MN?%�y�A�h6i8�C��l��TǙ0�j�u���!�@�'k�C&��K�*�`�fk���ԅ!�SH�fH���S�y(�jiA�4s�����jpc��f���I���L�w��65a��W'q���2i���ˌ�bZM���C�߃��ͬG��>�o�A#J-(؏�kjFUW[h���M}���^G"����5�\���cs8qt�V��<���k�O�}����IM��R��L�%|�Z&;Բd���n�L�&r��L�b�Ð�Gث�5 i ���l+u��m��Xb^��i�-;�����Ml�<�֗ϴm2�mu>��ƄZd���O���Ѷ+ڴU�׺�e��f٥�H{���SB=�n#�/C�R]L�0�؁�岱F����+��Ʒ���~���e�l*�]���8�u�𫄞�Q�:��Yjo2ۏ�^۔���A5.�,��pV��.+����T^�Y�M�0���-tN2Y(�0��r��
'M0Qֳۘ����UFS���j,�P��aY4�����dui�~і���V��ߚxdI���Θ�H:F?�}"�1FB��8S�U����)-ާn=��./���V���G�e��4Sd*�����O�{�g��NVN35����w�
K���"pH�,�7��i�A��	��H�`2Kx�KάAZO�DQ��*В�R�z�j�'�֮-#Z�E<�zS@�-��ż'�[� ������ �/��J3Rׁ�� ��C�@�H�z11[�"���-*b��h`��F�,�m�}��ɱ~�޸�'9�.�]>������u�X*�s��F�8�+>���N���;���ƫ�&fׄ%N�񥘇pR8\��LkU�R�he:�w������*>k{m����Y�O}�X�i�1�N2�1���ɵeT�u��n��:Hh�=�'%��BAu5�B�6O�P����&�[	�V�h�+&�Ә��Ѯ����db���_��6)x���v�%���.d�X=��NZ� D��D
�:�<s�3�IV��6N�"����vS�@����x�o"��[��񥅻�N�(8�`�!��)�^��4�k�i��7"04��3��˯<��~g�5���̛̂�i,
�b�n�jk�����8�L���w0A��60@���bv3+e��$$��w�bC
�5����:�`#��Z����`5�6F�OD4TX�BUD�X���>D�^2�5Ei�꾨1���)H0Ũ����4�T�txh���͑ڶ.i�Y�<�-��«3��A*���)��~ځ�T�"��LH���*D��(�XQW+ �)f.a"�)�[D��-)� ]�f(&b}4KQ��R٘���8/@a�5e3�X>-N����34�e�D5��aXn!sww(ҭ��#˜BVp�Vnx�r��U�K���`5)A2�׷���u�x,�����C!��|-G�ul��)�6��C��LB�1Z����c����������4_+y�`�3�
�;�u]I�
~6^�w�ąk:@3L�H�X��|L�c��J������Oy)=Y]n�1��Y�&�-��f<I���2X1E)J*����OBR= Z�R��,<�K%�4r�����|'�:k<��ӯ�i7bT���("��5D�Ю�3k�|��S�[�T0,�IBđa
ž*��3Q�[�#�N[���h�ֶN�K�Vw�X���`{�D
#���M����&�X��kGAZ8x��:�����CF���
b�"�6)�Ґ��'~䋞`�	���1²�nRL��<��w��
�rN;��W§@�%�b��W)�m>�`ȡR�J��!�wQItQS��sr?�k��j��o:�N:�q N�qau�l>1<Db�"�`'�$��t*JFY��z���̂y�@ik^"b�v�
@�:��M1K���KD�)���k�� HHp$
G�H�%��>	�l�LM���6H�ɺ2ӆyj����G� $��ќm�/�V�@���K����y	ݍ?����'��"��������9AI���T_��K�Aj'Ν������{�ރ�;��-�(�Kx�����e[qn~���}x��
�[�b�7m�B��£�/�#K��N+ ���xRqM� F�gK������N≓(�Q�D�$��vlB�kv1�gױ��i��SNۓ���G��9&s����9=��Ւ�� ��سic�Y�g�p��4h�ESI$Z�����"�i)��1�6`^GN��l�"tw�zp���M��$���38|4����݈�C�:>hCJ���C��p��Y,��.��v ޏ��Qcd6rX^^E�P!ΐ�V�ƾ�^C		g�f�7�/�j�2Ӊ�H�2���X�R�h���5�D�� �4��IG%��L'��L��pLL[�9��E?%%�m�%�N]�b."i��0]��5�/kH�,1[݋�i��:�Bр92Y!��z����
M,H��T��Pa<� ��>�#�$k�tb]��B�M������u�S�'񶫴�;�����T�?I�˯.P�5��GR1����9�gr���X$�	
/e-�j�l7��Ƣ$�xO�D��آ�b������hkr��ʊ_g۰���R.�Y��̽F>���A�l<B���D�����a#�1D/�i����#�7¤����T�ʈ&�.C�/��D�j	�v�1m�U�Sk+���2Nl&MS9��b�0@&5ڪ!A��+�pq.�c�$����c�����u1)�d)���6�01��6g�4�kS���P�Q`�8�T8���⌜��y'p	���G).���l��{��k7��q~tLP�����D��IPHyU ۦ��"��d�?]I����rmd)|�.f�P0ۼݳ������ti�4�l�<�����Oc]{#i�'��d~jw�B�Z�-�����49F�z����	鈏l��_?5.��8���23��@a孲�j^>�� f����<�f�V�D����%��؝��1ٔY1Ir�F����$� i(�B��:D<�RR?�6m�� Z:o��
�}/ݎ�������g>�O���YE*ż#!���(��?5�I
�@��r����mPk��+o؋M#C,���*�%�g���x��@ku�ւ:�%�7������s�x�4���n'lː�� R5�8і$�xq�+X�Pd�$����L�O���f��2��"�8�L���511�� S�����_j CK�1�m��X_M-=|����'����alD8A�E[�\�,����K�!�SW$�;	���-�G�V��k��bSSv#HN��sxM*)Z�%�O�}*x�u�6H�js6m���>
W8����SSE;��'�H%�8�Q2�8�}�@cu�,��ȹ<����D�=��΢�Ҽ0��A#����R6�V��^���T�B�*��#����E�BVz�7�(��1,���.N��w��*������B]h�@HLD����	k1�vam�S��E��FQ�W����^̵�g�E�5�i&��xc�&��C�
"�Μ��ǎ���U��A�m+KN���p>K�9�$���;�~S�I2���1
ug���sU��j�,.'C��4B�!��s��d��Az0n���*��z��JͭT^�]���uZ��!,K��?5
*0�Qsqnq�B�<htCA�A]�"~4�����y<x�A|��2򄜦�'�-�Ömנ�af>o��};0���J�|��8H!(�(�h���:�>��z4a��c��c�Sd�!2�ֆ�+��Ø�P+�!O�iܡ�m�����a��lB���A���'"򝘱�duk	3Ħ�U�	�饄��~q>2�YET��K��,���+ۂ�V����� �!�9�2:�(#%��v+�EeRY��6Q�Kx�1'�J[=fN!�S)xD�$�v��f&c|KےZ���D �>���$3j9L���V�Ǘ�s��%�K�'�I MQsL��++�Vi��l{�Odв�.��t;�b��E&����"װ
���3�ǊH 0���H �@%���/�(4�P�eH���ґ������X�Syg�����im[Ȁ��Ti�)�Mh%z���9J�
5WJU��x׵���7܈;7��g��� #�H0W�bc����*B�v�e�NL�z���"��vF����q�l���l3HQظ;�X-d���h�t�#H�A�O�r9���Q�pfF���f�T\+h��1��Q�c#�`�P"<��A�%E'=0�@�eh�z�PKK6�4�)���X�ր3S��R9Zh������o���)�mOO&]%���05"m2L�r%4�%���,,a�V%Lm� �p��19�z���K�E�N"��e&�h I����,�
xZ�.K6닎y�u(��[�*&���)ZLO3�X� S�����$�\1��8��Ѩ;���e�2��5jKR$\�R�)��&����\�,K����z+�zB�
$��R�O� ��J�P7f݉�|.3�PRBG_�~2��$+9��LC9Q�&C�}7�D��l
�����e/� ����ޭq�ػ��!��YG����ܘ����٬J*�@\g:	fJ�ĺ��,��o��۰�Q��R�rЄg�S����=YdV��f��8�NZ3Uݩ|�z��@r�Q}d�aJ|���@��HC����LL��iub��_��WK�ĿN���� ��059D�lcm��Z���P��I�/����{Z?d0��$��� *T2/,�Q�Ux�Kv��XIZ@�NgO/";��ݓml�A;��@`��!M!�Zc�4��#�@fY�q�Xp���E����C��dY5I+��H&N�'��s�b��H0+@��RIkǒx�1$=�L�a�x�\��,�/�$-ҥ�j�ώW "J�$)�9�Ѱ�x+oՀr��M`�Ru�K��v�I��Ӿn��:��vH�r��-u��d��U�`eW�Vgz>�j̥Vit�v|���;�Ɔ�N���i�$B>jE��-�	�iƛ����$�1tB	�	�d"��*�M�`Pk��*�TT9���m
!�d͠#0$tD��Ә<�I�*�A����T�gc���x�V&o�$���76P�j6�����n*�wް����P{&Se4ԙ���N:��G�@.���D���ĞQ����bϮ�X^��C���kw?l�r|�54�9�����4L�v��gC�00�mD�Evگ�XԘ5�h���B����fj�M��I�� 6o݁�͛1�F���gW�8��˳^�`}v	��
�A���k8��s�DzY�͓#��BD�
��0�dZ[1@Z�Oh~/�sE��e,-�Z:l9Cxi���0�y��&�w$�v�����e�鋚�
���㬫�G�tK@�U��	�T�&Lm��L\�gYr�H��F���Oh/.uqtPȔP�.�4E�����i�HmƎ�CԐ7��y����q��
��G'b�*�t�-�QГՒ� FL֍��_j���@|�tv)c:���q&f��]G������-*k '�L[���̚�]Y���O�]��c^�h;�G#R	X���7��՟ŵn�?|�+x��C�P�&�'�,ͯ"�����O�4�:��
Dq��j^�$^�r��Gn�����֗386��G��"�m���~+��R6(�H˴��-����%�?0�86Y��� fs-L�gY?*�1*0�:����
����#�?m��(�&7c<ՇZ-Kb��F�u��0��:^\���ŋ��yL6�p��Z�`a�mB�T]��7o�@j��@
���	�����svig�3�ֽ�fW���1:�.%bmX��y� �����.��5pE�ǋ�y|��*���r�2}1V/���0IJ�ڞ�5IF|�I�G��"�]F�>օ�v�㳎uW��M>Oex�Pšs)�����	9)8J���N��u�/�9i0]��G�d�A��{-���Z"	�Y�Y�Y���v����:�ZF��H*��4KI�,^�We1�Cߦ��я}���Ky|��vĴ�V �Ʃ�hs�l�LM����1�Μ�V�ڞ�7�k[��,\�u�A0���0Vr��4kF��$Q���M`�)м�n�2����Y�B
�T���C�e%����o��E�ֳ��7�K�F>5��kS[Y��R�����Y<qv���q�&���5<p�D��,V�P�/V�Xχ���>2��ؽ{+6�j������n��
#T���y�D���r���u>�� vp�86o�$�5 �F���`[��HD�V�mBk�BD[˫M�e��|�` ��m�b6O�b��	rÃ�DL֙��P*���QȘ�PmO}�5�Iع5��a$��������� ��c��5�����u�4�Lͧ^��j�*[�Z�'���ql� S���$�V�������Lal��0,�J.�4
Ԣ[^D�.Zm��	�������l�G߀�����<<��d��3[ȓ9jJ�C�$_��'܎��p��-x�+ @迮a[m�s��b��z�/A�ka��N)O�E+ˬ�i��	��!�Ch�RhRa�S�m���'�
�����wnZ���B�Fڪ�����>�a2���r˞ �Z��OS�����R�{Jx���sK�B�m��w܎_x��!��&|���1D�~�{"�� ��Je*K�6�̓�C�OS�����!\���㝷݌�v�B�T�<�
_���;/ٻ۩x$�!i��QduZl���=���u�6M�j���3��KZŞ�E��U�=��`ic��Bz#n�)��
�`���ٮS��ګ��T~���ba
�8aJ�%�b�w�Kq!��j���ڲz��7c��k�i���F�G���5�(�H��4SHD)`��b�X��-K(RI(gs�f�����@;74���ű3+x�L�3�f�QƣP�҆�to?���Gz'�k�Js4��Q��JX�����7�z/eۡ�ǡOт���֕'Ň�������I��w�(1o���MO����)/FT�j�!�(�mi�gX��P��(�%C^��\�h�4&�v�e ��n4l�V�b6�7c�0����qǱ����yT�`.�qZ�
y��o��3yJY_��1L&����v�BB;uOߺR��E�x�yIC1�ch���o��?D	2+��?Q�i�Ȩ�!��x3��LAJTmb�Ā�p���'�#-Ĵ~&�Lj���D@�7�C�Y�4ل� �t%�G�r���|���|3D�j�Kզmm�^�:Y*0"5WW
�4����I�d��8���9�� ��1DNW��\Vk74��<�5�k��q��<����M,��� ��ݟb|8�h,h[�*��j�"2*2׎��x6�Ŗ�c�PB�^��j��rזM�G#(ӂR�]��J�i}d��V��o ��μI#� i[�x1�"��!������+�v����b�r��k'����b��e��P�S(��v�D�߲s��i���*��� �2-	�8T�v�c߶��v�^��ʐ�����ս[��C��F�Q�X�<�8�]�M�,��⣛�s�����u	�|vS� &F�((t�@:�Sg��37	fO0w�-֫�W��Y�!��+���O��@��sՎt'ө+�U(��m�"�i��Ia��D���6���m	C�J������B�Íx�O�/��z;zJ�	gs9Z%Ό@�Wif���Ru�v�X\�����1�>ADSS�����mM������ē"�ڳ}q
F2�z~�N-�"��Y�$��:��o�!�Ww����	� �U"B+8�.&�H�����^�>���M+�A���r����О�#��F�Ғ��/棂�� ��:�7�|i�������D�\���'9�'1:�gV�v����@�C�WǂA���(7P,T����¥\89�3�����cj�0W��Y<|2���)�%��iԼi��e�����K>��>�ߦՋ�IH��93��$�;�y�عx�]�l0y�7�@/�+^���E|�Q��*Q��51y0����x�v~!ӱh&*��5:����'~)Q�(����g���W�!�h(��e�x5~k���t�`|�$��O@�u1�����0�\4�\k7P'�w(Z~
"m��*d��2(�����8�GסO�utV=�Ґ�f\6J��N$h�SSk!�je~Ơ��$�H0����"�5�;��x��8y�k��X����y"#�l��[�B���= �l�Z�^������U8aC�w��2]�[;-i���/�iٚ�l���q�J��E�14��.]���4j�E���y˘�,9�O��eE�S���p�hm���8�2jc�(�����)l�699:HfE2��(���}H��j7���O����R�K���.�@Z�#�2���9,-^��]B4���d4�!
��f���cv�]GL���z6�Vj�nm�D͗�Iq}��
�Xݖn�	 p!����skT��Pغ��4�����F��^ƞ�A��`9��ё�d��0p*Hk�<�Vo�0H҂��36�����}���FסT��>�~
Mc Ծ��8a �.k"���8a[	��X(b��%�ц�||p C�Y�����b;�	O�?� �g������1� ��p�W�*���)�(&Ȝ�",;��4&������VZLC��-š���qSi�h��d>,c�<Vxi�n�a8��=�8�Z\ 3uNL-�2�=6ޗĞ�죟"~�Liަ�d�'�4��-��75�����`hl�ʪ!��	a2G-����#:l�fuB,#��H
��0�֖[���0@\ڳe�^�;����'�S�S�så�8q^0�r���r5�����<-��J {�(L�S�tcr8�TPEm+�&�E����WO2jg1�3�����"�ur��X2̲�Ր)�0�����<�����7�x_}dw/�k���E7�:�]�iΧ�k����$ܢ� -`_m)>-te;�hGm�6�O�^��#tԀ�sl�g�I�H������#��o�ye��Oō�����s�$(,��1[�o��P=M��JGάB�>k�8y�_��;�J��t9���|$L��8�W�˷*��Y�+�BYH�'?q�,���"2
���%g�Ȫ>z;��ց�.�����0Z�'�ݸ�8�d<-��ԅzyj��j�myJGu?[U�
*Ԧ��a�{�Z�L=���5z�z�J>J�P�����hG;US[�ju���aV4��V����:�F�,�����:+)Ӝ�����9
��0��͢��M3���.K����v*��l-�]��ڀ�V�	�j`�&�����'�K����N���K����#��c��8�^���)MFK&�c�0�M|L�A�l���T���e~12�~
i����5A�yn2!��&��I��&���R��� �"12l�j]�d����A��H�"���M��e0��4oh�\�� @K���u�_�����y�+��m[��>�H� *�"L�>DMK������MkG۱�t�q�G��w�\�G���I��<��p��=Â��DU0�p��Ӵ}/-�|~ٕE��:���DLV���P�Au����8A�|�4Y>j[a�����}�6�P"����<!
���x̍�#dd��� ߇�)H�WS��0z27�#��	.M���FnE��?4Wd���aK�$��ߘ8�/�A!�M+ʦi^Ҭ����m]�+�@�C�x]Z_�3��ƹ�����SX���ųgp��i,M_���j{/R1�vl�.Z/�L�Hc;��x<B�0�?��� �M�J�C�#��PH��u���U4���xi��}����&ǆl�F��e];���O��"e۱����iK_4�0r��ŝ���6E�Ck_K'���P:��{vc����l$���uL�����j��a�G�&)t��� �Q�n�4A��ap8���1���w̿�� �R��\��*j���u
R��m���Қ�ޡŊ-y���x��wC��<S��f��K�Q�ґr�(��s%�6fΟ��ؑ5�/&�	T:bD8��P�`����B��^c26�M�-���v���]�t��3J�e�z���L���н�2!�8*�)�/���|�ׂ~��	��9�3|ϳ9	zip"�j�����/�JSi�EM��%s�e�.��������\S�!Ӕ���3�2:��\�Eg��C�I���}��a�{zr�r�9ǽ�{�Xb�II)Z�,��l�l�˥rY®�����U6-�d��D$�	"�����ݛs�r��or����n�~�鹻�m����y�	�y��{µܸ���ݹ�[Wcp�jT�܍
q��M�_��q�|��|7?z'�y������z7���Ť��x%�޻��~L�0��8:|ݏ�F��_���"��w��`��e���J�n8E6>�*�r趍��r��6��+/���B�FW0�A��(X���Qp	A�px�#%Oܔ������0����y,��q�YXcM@�y�T+�%��P������T��i� �;�����+3��(4��M�}�'��f����Q�G�kцQ.�n��_^l��^�L#�G�'��%�Ц0P�2�g��=Uvi��}�,C "��fQ��s���·�AU<3��,��ݷ�k����Y/�{�������x�ᇣyj9����:�g�%<��o�4)M��jM^�B�A5���a����(*�iq~	�/�ݜE�f1,P65�ҡ���OA�Spv�����&w��&B�5�(�I�4���U���(�O��\��N���ޮ�k��[�8t򀌬B���6�G[��/WM��.��j#��2S%�'5B�h'��ˆ�R!D�ǝZl�G����������+����}�n�Ż������މ�:�{��ozR(s=c���l4PK0qΐ��[Ӵ�J������Nǹ��4\�ϝ�������.�����ݻq�����P�ư�G�=�E?	"��*Կ|+Qi(9�KgC��ho;v0.�X��=;Y�&m679�3�q��\�����RL�z?��H�G�t3�w�������].	0�蘸�ȭ^�P��iϞA�P�����U�-�~��(��7Lp6��a�#Bz8�iH/A�뚁��K8�"��z8+�U9Y�ۏ���8�"��
�xG��g�˥kN�x���+ή4�.�^K��,����3�\�wq�{�K�T�N��<T4��?�d	v5��+ܤU�^$t?:N ��/����V�W��� $L )�@�� ��սۏ��N�n/*�n4���}���������߈�[��n�������]�x'[1�9���q,R�Y���#�6!�����b�ڋ�V?���l��=��ɰ���~X���ݘ���A/��QE46(a��9����0���:.8*�L� i
���d?�y e�`g�@"�A����(�a����F�j���ǆ��=؂�`"P���:L4ߞ��/ǅs����P3�xlbX�2ĺ�������B��Q:��������sS�X:��N�#\�E��EQ�oa u�Ӌ�*�v���fט��l���oo"`�1���!T#.���y,�]x0��w�3�4DXH�= r��j���mMbeBpβ����<�Yх��

Y���N��&b�94��G��^'VQ�Nb�l�"<�����X9��{���4�E���T2y���o���@�\�}+���.��~�Pl��9�֝6ۓ5��L,�I[��Vn+᎖��c/Gn���[�@x��$qG���ۜ7�(��&i���!7IC�JC��60Jr9
,$m�*�uL%.���+�'�0I[ԙԓ:�O�DC;Ԫv���k�t>*�½����ugA���Pv��d�~��?��{�X��[X�����I<V�
N��kٮp�|x��Ϟ���0�W:�Kx ��?x(���\6 x���K
c{s3�~�I��Y���%����ʩ�x����C��G�����[���w� 9��z���Jf�s2���ю���*�����.����X��}��[(i���|Z��`5�a��!�Ĺ�y��v.��
�q퓛ػw�s�mcgN͡Xgh.����g�u��L����`4��:���K!����Ae���� ��=����2���ݡ��Vc��B�G�..�@a���K���N��a�߲]�
�bi(�iQ���_D�_�(w��q��W�\��R1�?i��p�4W����1N~��^%Y���L�}z\��P�jz,��eΐ�Wz`�m��Of�~�-��`4��kFt��~T�a�Z/n�*tm�%;��n�<�����{EM��w `wv��QVn��6��o��·:*�� ˫�V�眛�����sp}�9��u<-⌀a�(Z�`ܣ��-,Z`��X�|G��Z[������pɐ*�!��cf-c��d�T��"�VC��b6�e�`������>�p����o�a+6��bsk-�f�����≧����{2Z�eR���m��^`��*�Auog�X�X��}����ٍ���8�l���q���1������nj: �bRI��;x�7o]�-�g��"���x����Pb��������1��=:D���!*&u�MG��u��
�s������P&  dzwj�#$�varn9�x����ch�.'��\�|�.����o7�� ���#k�i��Θ��(�w�����q�9a�.x�U��x?Ϝ���Ӕ� � 5�;A,�2@@�q�w�ׯ]-]T������ZG��KrC�*�]/���v��}�B�M؀ˍ���-MXa�B�}�VL�9
J��F��۟o\��l_ �q6y���@�����s����X�����w+(���/a���M�#����^x%��jC{X�zhy�C>wn\����ՕX��a�LUcq/��w��vEyrv#�j�>��̥
��m167o����{W>��x�n�����#��.�g�~4�|�B����C�����.�u��c�+���B+4�Gv�b4mc���������Q��Gב��F��nlčk�G��N�މ�~x%�]�W����ۛ��J����^�\zJ��c��q�G�FCʝVSҮC�a�-<.�Y~KV���wG��ެ|���d8_r����k������]�.4;�̽�"H�#�A2A'�V��B�����HH&9?���v�&UY�xYFF��r�<aV�Y���8*��!���\��
(�*kK�o��������[;����8�AJI;D�['5<Bܥo\�����İ҉����O]��zt9���g��뛱�֭�n`=߽	���-19�F��ƨ�P��y�z(��xr��Ou�
��T���4X�9r1��:p:h\WF����vh�:�8W�m���݊*ֹ�߭��zT��Q;�, A!b$P��������)da༃����UIc]ձ��vfa:Vo�Ǎw���Z������D��
=�|o}?n��d�{��Z�o
�\B���̮л�}��G�R�z1��x2x�nI�E�C<��p&�Q��N������B}���c�x;��������a�r�Ɲ�ygX���m,Q�B�B��p��m"��m=��(����9D!�x6 ���N���Mk.����<�M�]����q5��u<�V�\��^�^ߨ҈k�vcso"��6�f�ü
�Jl���¾7����7̜��ۼA����Ҿ;�uc};:�u����m�%���>��Vܸ���T�k�x����r^����+(��E��H���Fģ�Z�p
U�V�ɘ�d6���2I!�2���yv���PHz2�����r�/�e^��0<����E���J��H&��>v��W�ۚLa����u����c��ͅsi$��P����wV��ߊ�^{?�V��7cum-�7�c���m��k����Wcm��Nۓ�ǣ(�;=���06���Wo����Ц�v�=�^���n\�r;�pۍ)GJ�9��>�K��������x����[W���n�DV��w��[�qonT��N��k���;>�Ro�Km�w�W�6s��7�Ïo��׷�;�qs��唠�յ-pOӖ;;]�jo��i;�BlP�n�!��3���D�Y
�T�pZ�*� ���à��a���Uk���z�]G��S�٪�����-J­N�W��=�UT<�3�R¸l����>�0 �t�J�:�Ðr����ݔ0��
�zr��xҤe�h8�X���(Y�	�c��K2O�9��*��p�k�ފ���{�	��>$c�Zi(P�ZG�5�頿��/�RܿP�-��X����_��ˈ���%lDe��� ���b�>�3�(V 9��׀µ�)���q�|#.O��������bU�da?�Ri�l�)�T�w!�+WW�S͘�?Cj�������m`s���.�@
[e#"�zr�L�Ħ p�+7h18h��#�-�G�Vc��{E�@����x��t���0�����C99��}�g��ўo�w���ql�;�;{1?�;�<%�)nf�����E?<;j�V�]i��������4�|����nT���]�&,H��3�x��"^=��)��(gkOB�� �(�����ukz� �N8JF�:k"�g[1�O��c���w����s�j� �=t�f�j�<ܗ��[��Of��G�l�8�|�(����sX���Rh� ��m�6�Hуڧ�{s.
q���mm�f1���Sj���PR�{X�ۛn�7��Chw��X��E�_G��͕.�ݭn`�U.��4��Bs��N�������s�8E�V�2�٨.COx�<Ml��xG�6�*�U����e6�%��O�~
�θ�s>��D�R	��]��CXX�~�� �a�z��k?�|�}�,FV�ݶ�����b��)ol���F��
���xK�+�=7��܊��a�c�-���ѡ�D nubmu!��G���q�\m�/ZMh�Q�F�V��(G�t�q�s�m��\#�A=�c�2Wi�q��L�w߹8��?FA��N��N x�0��q�ѽ͸��䁀>��c+-��^.4���;]�������hw�x���{F����_�����ع���>w6>���l,��;���%p�օ�P>(���j�
��s�RY��x�+I+��Qл��x�K�A�L$����x@]�;�'G���ݒ�O����|�w"���ݦ��#iL��N�=4zQ� AKҪ+�;�V�"��䫊��(ڠ�s�>��Ŋs'e#h#����x{���k 2y�}=jL�6�Hy�q�{����?|k5������==W8��
4���*GN�����+gb7�O���q�&�51Wwo�����z��x�b�9�W��eo��f�s�z����� ��Ҧ��5�@�ن-�?�����x쾅x�W���_������ ���������Sq���X\:�B�o���om����fi9jg�� /�9}�'����}�n��c D�������O��t-�c "pQΣ��~Lksf2�'��y�a���},�lZ�����F������޽��!\��!�0�r5h�'�ޡ}� �]
:��
!d�;�U��3��;�Љx�8��\g�p����s���N�nC�k�E�	��>lw�uֵDf'��PlZ�x` ���j�W��Q�5�%���U����3m�^'z���I���U��¯<�X'��I�*�ý�t��YRq}�h2QxW�~������ǇW�c�.i)�?��d�L��^~��=���za�|�d�r����M\�m��NY8JO�3���W�ڏ���̎�c���7prVH(��!#�#��g�V�G%�#�2£�+
h�l��P���٨,;�z�(ND���h�����7;$-�w
��;y$"��T�.EP�\�w�TN����B�`QĚ��`OF֓r�-�F&���
�(�x�#�)l�}(4z�vD��v�bP�3Q;==Hϭ\����>~Q�A�9q|m=F�\G��H�2W*b��^�m�Y�H�]�*�p���`U7�bp�vT���>���
krc��J�^���b�W�L�!��+Nl �	(�mK=���A�,uU\5�&��(A?<\�%�����k��9`d��g��#�l7�����99�௔L��K Ic:�h[=sIA����� ��P���&�U��A|�r�s�ϰG3�zo�ro������v�~�pȹ;Ӥ�11�Th�;2
����F{��ݷ>�C��T�3(��?D��B�:W�_|�x���q�`t��㹧/�?+�^�/>�H<u�x����_��B���?�5�q�}���ع-��j܊Xì% �8������k��g�~@����k�5���}��gf� �g�}6.^�o����q�ӱ�0����w'-e@�\����%O�]a!��]$�p N�ψjC"��6�ݏ��VPh@ �M�o����}W��+���+������r����M�La��5r��J�o|�K'I�Ǚ��~P��}vT���c�n]�����KK�<�})w�11�=@X9a�CK�:��_�Hz�_��_�>��Zddmw�g��o�~�w8p��	ϛ�:ʾ�v�X�Ʉ~�A1�1&ړ����P5�Md�*<���顈w�l�]K�2ް� �A�I�{�������(C*.���(��ȏ��N�N^���b<�j�@�D�mp�) a���rg�|m���!�7�[����fKˀgۢ:".ߙ��OE�Tr���'��U4�2�	u�I��ѧ�0@H�i",%T������� s0	�#�h�By�t�A*/�Z�P�;�%�5I��,�sJ�Q���6�R��/s�Q[���B�Z�ٶ��X���+�sG�W�t
�~�GL=��:�7W�GPe�@H�d�oh7��c����Lph��^ȡ�+�9<_\��� Ǫ*B=!\=���{�َ���9 �z�"m/H~�3�m�m\�@ Oړ24��T*.R���+�k�h'�Wߏ��W1?J�<1�����E�)��
��5yMZP�kC|�����ɑ�O�*.�:�ٖ[���ҀZE}�E q��d)/o�C=5\,�|�����G$�8�"�a�2M��*J��(��N���|�����l$��aW�>������O?�<�p|�g�g��j��K/�W>���ڗ�/��b<����ckw��F���kqw�7 ��o
壽�RI��f���G�Ƴ\�a�ͷ���;[;�?�S���Gq9iP�qy��L�+��wo��YkR�����K����O��Z��g@>@��S_�q����bQ��r�qq>�{�4d�a>(���k(=-�8�/[��!�~�u��	���������(W�U�����h$�A�K�\���*�FFM���#|�m��]�U&`Zʭ9�|n
���yᄨmV�?�4%��c� ,�.ʴ�Ck_�����٢�*�O?��=�QI?Z�X��U%�s'-�9����6
�5��ZG��E��+�<�؛�( �5<���SSѤ�!�c��p$~��S�A�.f�L�I�.p8L�zW�����84'x��.SX��Y&�-�w!E0d^Я�FښKNM#�f�b���]�*�!�@'2.xWP���l]G����3 s�`ާ�m����0��"ַrM�R��t\/LgwU�b�(T+%WۮJ6<����`?8�'�1u�����9Կ��uO([告��9G陿ߑ��F��bzz6Zо�;�O����m�v��Q[�E�@��Q����B��i����Ũp�����|@й��"�0j�d��<���1��5A��	pU����iۺs�(ڟ�]\�z�z�*W��),Q��D�"+��NvQdy!0������XnW	��t1�2�)��͐ԅ�)w�si����W��y�`=��cf�<�v �="��yy��٧f���Kr9�䆃(��|ϥ���^�mS��x�Q�����K��#�hC;p��������|o��zƓ�>=�T�	O���k�7�/��P2��1�� �`?�Am��=��Q���������?�k_AI�ԙ�(��&Z �`駠��ߋo�������?�o��j��s*��D� r���ͅ���K���^|4^z�r,O⽷ވ��Jܼ{��2�z�����e�q��3g�@������W?�k{3qP=��.D��Y,۩�͎��n��ǽ ;�#7C!§��q~����ʨD��ۉ�Νp?b?�̨6����z����GU�+�׎�9���8+xu������rm��MrGJ�?@1:�JjO))�"��٫�`v�̑^���%ܹ�8¥���������8�7˦\��x�������SZ-<r��C�����Q�6('WH�6�?�d-&<��H#N<�;����99�nH���^A�u�;@��k¯��$�܋!� O��PK�tM�߂�t����H<��H3�9w(��U�B8�z�[-m^�K�D��(e���0oR�Y��n�|g��CϞ�'��~Z�❺��k��@uQ���;6{��4��qi>`����mӾ���u�+g�r��T��� bc-F^I�r�%����������sg#��kh�^
��GG��݉�G��gpc)IK �0^��4-5Pb��hei^�]+)Yz�+8幼A���?	>�c;���r/�.|�q������HZ�Q���+����Z[�S���|t��z ��
�%0���>���vTo��@�w�9�zz�u��
�f�)�r1Nj�ˀ ��b�G1��Nt�il<��1��2�ȑ���<m��kV�f���(]G4�������XYl�N��ލ�k���LΠ5^��n78!�UЁ=5��x'j����J��g�y橸�ۊ����ʕZRa���m�|9�@�@��6��� �罋�|��״)�ElD�q!޲�\)C��se�Գ�`��t* �C1�({���{��	Y!��la�t����9����F(�~��w���[=?#�
��8��� ������η��^��^�G8��Ր � '!�x?`�o^�{w����w~�?�?z������9�a״�֘Y9Rk�y��s�����م��wc�{w5�vV�ϱ�:�E�gk�0�w�X9�,�y}��r�k�r���0��,0Y��*S�C
!�<s��Fc�v3x�x{�v�R����� �n�k��В�0	x2
D�Up�v�-g��Ff����b%��ൡh|U" ���ՕT>I
.���0�n�CeO�9���z�v<~�cI��Bę��a�;��]]=|�t<��M��i���%:7��FezʱUٯ,�:��5�$&?��uJ&��\ਟ��5r]*=n� �*����}�!Fƞ6Jb�ò߸����by:��9@�c�?��5��n�M�s�C_eE|���u�ﭫrW�w�U3��d�(M-w�p�W�a�2G�8�46���=��n�+�F�q�~�Z@$�	{�ʵMi���MeeԱp�e�N�e߻s|�"z�(��\��;� ��"��<b)x��sQ}���-(1xh���T8\���:­���#�HQz����T��[��p��OVڢ���*&@$����tO��I�*�t؁����rt�舠,�Z�g� �6�z*�{��Ƽݝ��!^e�37��ů�%�@��"�gض�[kQ�~��:�~06�v��/Et0��@:G���[l�8�%�|�y��ǠJ�W�7�>rι�~SRi,�>��ףND���Юhi4�㹋���9ǳn|������N�ަ���R�jx�8U�#�ܢ|�Y
Z4f�ho¿wS!_��X4���Gqw_#zS.@���Q4'���W�����S�>�&bC�!�1*i^���e4��M���/�O�I�^��'y�^,4k�3p?��M��d6<_�b�F۶��Y��︎�3�dF�%�k+��,( �Js�	2+�g>s>.�u�`{=5:ՠ �(���ZpZ��X�a7|�h�[��o~76�����ݨ�
-�h���Aİ9���j����D��n�c��t��\<��C9O�%�[S��5�՝����7���V���Y����!��A�!��'y0+M�iU��\�=���V�"X�� �a|M#1θ��J�)��.{�=�b�%�:��u�&������T�J��\���F��3�lW� f3T-���&n�k�kMe�Jc���1��2k���qp0�3�97}������(3ς�3����)�Բ��z;�@�8���k?y Ԇ�]`�������U"�m=�u����c�� q �Ch�=����N�E8��O�W^z&�;���/V~,z��8 ��П�#2��%b�ekv��=Bp��]Anv��D*�?F�Ԁo�`�|L]�z�xa���b�:�A�}'�]D`���*�Oldp ���A�#�@�ܥ23�A>�H�G`����}.���\q[���2���t΋]�y�r��(��B�Y�:mb �����[qz����"�]7\`
���ȩ�"TƗ�)��6��x}�Q��sB� �Ih	��4\�C���k��K�k�'��:L��PG�wb�s-�G�P�������A]U
U��_���"k�V-��M��j�`)��M@OYf�</W�j���� �4�5	S)��v�ANC��`e��
�:b��wHp?��W��%�[ ��򠘜 �37L��1D����cy�o��A���X�(͉����UR�<�G:А�"��iI�\�q�����.c >��ӱ�_�����p$�$��W�O��r�:�|�x�,mZ|9�mDwڄT�=M��\[�2z��ˡ���0Kn�ķ��:�a��W�w�OZ���JD�Q�)w� O ����ˑZ��%c���60�w��w��g�>�pZ�N;�W�܋?����]��^ܾu�8�q��v�k����p�:���Z8�jW�Z�תnNN�,x��CآأX��ǥ�������/�Ή����;�ep�{��cc�NA�����-���Z(�������ßm`��~�X��F�����:u�����}�I�u�D
��}��{�����d�Ց{��q�*�N����M^�.�F"(\�C��p��Y .M8"���GXpEpP�]�o����Db�B�i�S3�S9۾6��Ǧ�x��Q\����j��ZF!؝�b�v��\oÉq=�ӎS8S�� a=��d8���s�G�)`C�7�[1�4��/����N��()Lz0~*CD�f�� 62˶�� L��73w_��x� ,��S�a�]
�u��ֻ?��B����r�r��4��8l�\F$���y*q�s`���ԁ�ļB�+��G��	�V�R&���Yz���+(���v\�)Οj�b��$|R��q�V�W�����V���}+M�f>�N!�{d����hQ�T-C.HE���������x���#�H� �A�Q~�ʿ��Ԫ�b�=�%�)�,א#8���7�*��V�K�Z���h����W\"��;�^�� "�`�O@ܹ�R�0-��~�:��4n��y�L�^�	r��<)]��𝆈��:W,���ٴ��$0-���V&��sӱ��o�،�n�r�'�RX���T������M�{���nu1�&���ĥ��׎kk����2���U��z7�L!$L���\Y�|����{��}a_�YJ���(����34~��MČ�	�<�q၌���*��xU������x��^����`�� u�+���%���� ��ӟ]��񗟍�.��(S�������n�ŋO?�3�qzy9f������x��/�j�F>��ߗ�m��N�g���<V��K��3�8�7s���8�-��bei)����X^\��g�����Nl��Ɲ�8<8"����&ff�<�o,��b�{�x:E��mGk��S��I��Q��^�$���bu-d�"P�+�r0c�àKz	�3:�|���gy=�~��	:R,�g;2!4Ra�BTAAp��.w��>q��̟�#z;ݨtbR��>@�M���r���� ���!�{Q;<���xl͘��ѫd|�̛�*)8��`��K(M
��K�v'�c	/�C�*>��u��e^w�;j�k� v����`2��6���T�ٽ�r#?�kj�Y��<����N�Q��&=j���CK
Ө@E����2I։c���ΐ�w�2����'e+�j�1Ù�
��Ł���%��%�K��;'�ʯ�F�ra� *w7I�5?�ٕ�x�KO�Xܽ�Nlch]�z5�?��}'�{�1ܼ���8?W��=u|�+/��s�u���qA��ܘ�Þ�E��%��^O<@� ��]Yg�{i��G���y���G\�3*�fHU�08���:G�9� œ�H}G5j��񜧖�G
X�OI_ƧLۙ��%�9�6�<�����l���1�x\'m���/���Ao}?����{�Vi����c96�@��� @⿇E�@���z�����3s������8L�^c��(��hZw֡�~TE	Kҝ���XC7w6�uE���ڭ/���@S�g��23�Wpaқ��l8�Q���L��p���eÎ�8UD��;3_&�c\�}����z�g}l�=G�ꢊ���a1�o��F��[E���7�cl"KvYm4�j#>�A kgb5a�wn��:�g��.;�!��X�`�z	#��?�Q��	�m,�p����O�d�<v!^|��x��'��۹++3x<�q��R<������>�����k��s������&⻽�w�Ć�|�S/:B�M	�,��RI��[���#h��,��GͽW��b�J��Tb'
�RA\��������0��G���ZUv�9|�b�(uW	�@K%=�
�
����JK�u����|s�$�F��JˠI��7Q$vS)��iZ�>�Nmu�u��qgX�(��j����{�
8�,ŊyA<�'�Ju���*@�N����P�-��Cg<��ߍ[kGqg�ۛ�qx�N�z��X��1?1D�@���O1��
�Y`'ne�Tm��]x҇��,*�:�#�(ۙ�!=�dN����՜�m0��̐�,i��e�<x�S����8mv�%]�9tV<Vډs���N3�� ��#�:�LZn���\+~�'�?�3/��|���;�>���'q��qLwo���kQY}+zw?���F���1Y;��<u..�Ǡs�>�� >p@����ihL�kb�f���{�*+������ݖ􌐗w��d5Gx ����Wr��Aמ�yho�:a)�	)�mC�N��<̟r)Gb�>��?L�O���6��T�G�S���JU�8���� q�݈�wc��Iw�A�hC���T�R���y�ҩ�&�:N�M�ŕv������X�Q'��x�s�#��U�k+��*&����}0Ys�����('��]�%���3��_Q�ރ{�T%��IR_���{�(7��~���	]�Q�4M	b0����9��r��qr����������u���ܸ�Z8W~XGx��0�\
GW\e��+4�m��
�~{x/6�.��G��x&>��������Ʒ�î��{�ڭ�B3�>���Ppتk�AU�v=.<r&>��C��?��?�3�W���W�+���O�J�3�՘kUcv�͸xv�h�g2N��N���� ?2�PS>���Ƅ�jP�����B��87C�캪�h�fT6*�Eeؤ�!=#p��M�C^*����Ŀ:��}�i��a���+#C�Z���Z�}��]k�J�lgw]E]��|�z�e�b�ܫ�=B��s
S�Dq(����~b��6h���\��i�$����w���6Ԛ�٠����Ϯ2Δg���x5$Ǥ�O�n�w.;����|���B����x���8[���H�c͔R��^�ŘQ�X3�&|E�X��r�e�%,<ˑ�<O�_�{��B�4㐞��'���)k�2�]v��;��'��;J�
�R�X�RD!��@�Qs޶J�{��O}L�����SX�����/ė��x,�'���^�Q�噅��W_���7�l<��Ř_:��pW��X�s/�~����+��M<Kw��]oX� TN�;�w*���N��wP��.Д�3��y^�M�]o��N� ި淣�Q�{<��˱_Ce��uG�C���PO��<��a��Ͳ�N�����s��]䜫)�up
���I�� 3I>���~�ߏ�g�#V��qq�z������i��v(�߃�i&�'��{�����][��8`���F��H%>y�q`U�e����Cq]A��֓v��nT$N�ȹP�tiOE�b�}龤J�˷���X��*i���`n��s�#N�g���ó)��'��wR��.��s�9���~\���ɳ|�c�N�cF*��N2�!����G �����^�������k�H�*&�8}���>@pFs��+��g�C���Vm�b��l<���x�X²�i:����ٍ��z�mrފ��Fr�}vo��d�����؝du(c��v�A!D�������MKG���o!�	����ri��X9!K�$rM.��Yfu�����n�"nS����֣�v�N�w����VN[l���� z�w��y��t��;��Gnu��D�ԚP�#�tˏP�G.J&3&����TYgaX	8�ߜ���X�p�f��L.I�&���OF�Q�e�y��9��d͘�I�����-�����x��r<|j:��w�.m8Ʊ]���C��P����e���T �
IᖔF����3�>�QOO\[G�m �T��O<�^���=�(D��	�Np�x�
($����uz����Z[7��Ғ�:�Q�[�"}�Ω�ti9Ο?ܸ�#�Vf����c��r�{����K137E�Z|ts/^y�j|��u��8���BV&�{d1Pl\k+�����S=�ԩ�5`LQOG�6�����\���:ʕ �{�(
踶���8���D�9oK>өY8H)=�>K� t'����&��FE:�^@�o�E=S�����+���4J�-Nfg�9��i�0I�9Ljҥ�J:�&�陑��
?[�f'n �m,�Psr<eϬ����o�%Hc�_��lsQ�g�&�5�rn�
��_�%9䧀q�'|`K���S�mdM�-1�'���X��������cG* 2�Ѡ��4啁��a�LӉ��Oy����!a�L��C�Da�`��4Z��<�G�y�x��TL!�G�x�h�Uی��XވݸJʻ g��+!_'�O��Ӡ�XA���������9ӎ����t3n�;�m���;�~-V����j��W���^���+��ۯ�[o�0���{o��w�DG
q�A"�) #���#��PF���p��M�L�G�ݿݍw�{��wV��2rQQ�"I�R��l�ޤ��(W'�6`�%YȠ���@頀��V�s����~5�� Y�!���L�.>;:R�@X
s����E鮾������a�:�Id�������r�=0YW6��JT6�i�8�?�z�{�J""��æOS��dH�S �L~�sG�T:����K�|����(��nM���LL��1~f��X��$y7��\mE�>�Gոӡx��4�pp$c���P��`���:>Q>�[�q�ԛ�`M%J��$X��(,h'����EN]m�j�\p��6���+3/�ϠpT�XNQf9�?��*g�[�szW�<��a>I�\+�����9Y�٬���aܾ��汾'�s�ba~8��OǗ�/����_����X�p��ǽn-Z�����<O?�x�=�HN�P hB�+[�n�c��A������a4p�\�	0��h�����Q�>�������������@�R��,��E�	�#��*�$�BOc�4�_@ �lI�Ȓ��m^��nvge70���<��UXM���%��LO���}�i=+k �dE��D��;���JH��~^6ɕ{{��O�ŕU{�0�+в�2I��^XWmN�Mإ+h�Y�`�+?���4��\�c�Ai�^Kg�,�4ϴY GF���y�N	�޺�3ҧ��NT��_pu��cEΥw%���"���x>�r|�������.�վ��_�����{�|]
�a!�dW�>D�T���/<��N�8��I|���I�~\ى��Q̢��y������ƾ��G�~���a�)>�S�1{n>.?x&�0ԇ�H�'���98��[��������?�n�����z������ko����z|��?���Zl�����lܹ��V�HK1�v�f��@hO!�]���3���aR #|��Do;�7?BA���5,��Xo�e]))���n���&�%@@��V��J�~����@nE�����8���?��9��	q���6�gc��!�_Aix����u�D��s(煅�h�,ƞ]9P���j!� ,��l�쪒�i�a��m��4G�������9�g/�x��_s+������i��J�
P��F�,�����_
'o�J�{˚�=�J	S�d�B�>k���㒞���93=�f�PB[G��:0~a�q���p�>e:�RQ 0
[�oJbB��LϽ�^8��] �T�6���I��0��lv�y/�1�7J�@����I��.���#��;�v7���CAcx�_�$�!_=l��v)�o���k�O,Nţ�brr��<��8�&x���X9{&旗b_³�\��
ʾ�qxwo/'#_�K��m��ތkW������f�7
����ս���>T��x�H�pm�Gs�P��Q�d�V*/`癫H+6�J$�m����(��ھ����h��B��}g�1h��[�������#��t4��/n��55?�]��B;��q�u�P� m��ʫZ��6�p0G�M�C3�f�Vh@� ���И@`%�ٻ�vx�wz���]�3BE1�-�ܟЙJͧ�WAH^���L^ �
GZ�mү�CL'}��rO�ä�-�3���,��r�&7i�_j��l�����Rc�����"�v#79p��E�Ũ{����U!j��B���b,�<�_18���o|�����W������#2h����a��b��F��O?�F'zd숤V�.���΅�|�Ѡ1���K�!��^y��������@���,x>f.N�C�����||�sk�b
��P����V����w��z9������ׯǫ܈�?�ocu�wu3�������ʍ��r������F76�hRjT�QuT��l*ޏ�.�y,�v��ɜ[Њ�v�Dm�V�L<���ݛ��\��Qo^�«�S��la��益����M��Ǉ��Q9�s�4VkFy�tK�J�EB��d�������O/5���s�=w&|�Ѩ�����!��(<���L���h%�T0�L}L���L�MKǅ�v������7X'nmn&��H0ٕ� ��uL�VX��$v�72��*���
���gnIƵp�h�tGq� ���N��|$G�=�$uN�'d�L����㤛&�
�!��eC>�\��b��L��K�r>Ik]¬'��<̛�K�%�����76b�/��'�9�e�f�6�ē�8�<n�z.��)p�+|v͐k/�]���FT���)<I}�Al�ߎg�x8{��8s�\�̶cfzzi�d�S�Y�u��b��p�q�F|����@+ҶU<��k�U����Z��o[���Е/�-U�w�?��i,�������1��D���bދ�+ߑmzI~����Zg �;�8�.����#�ո-�:A"o[� \ǛN�š<���X���n�Y�!�=�^Q`�-������sΒ���C�x�����^���V!i�8��൧�^j�p�^R�W�M��%m2)�H"+뒼t�`nf����Yy
�����5��HE�������I��ۥEW>/�%6����w��=>�CZ.��i�#Ss�$���ՠ��:(KR�x4bˤ{*T�����Q��2M�B��?ڠ�q|��l���?1;/-���N>�8�H��ʣ��+�ߨ���h��l��C�X��F, �"�9_� ��c/dazi�؊�;����	?�#8<�ُﾳǭ���~&���>�|�y�9��B��}�/�d\�|��k�UP�����d�]/L4���B�y%�]7(�� �	'tN�`aΜB9.� $�I��7�ՠ
e=�usul��%\d���!R� ��a���R.Fcz%Z���VN���f`N��n~?p���-��٘�B��VH�?�vjj�y�p٩[v��'m��\?,W����\�gY�V+m�nI$?P�R��ϧ�K��q�Ae-����I]y�������VhyX{�����.ۣ �A���9YPXJ�9s.p�p�2�x�+�:�C�%<��a���i�gY�.�E��Oo�A8ʽ�6H@��l��x.�P�� ��4��FGQ;ZGh���kqvz+&��E���09�#�1S�?e~δO�1��<y���#�{6}�BN�=�0KK3(�8=��.��g�/�����3�?��Sq��z�޼A^~t쿦OM���X� ���l���P8��t��/i�a�ҋx��iql�� }�j�m��գ#�����\R+�(�s��^�؎�6����4b�:�|���6�\�SO7��3咟���r�
���b���z+n���H:Ѩ�"���T~.a.p��3�g���|,6��
�?꾒N-K��k�d��rN���2X��B���	��*qf�<��)���b (+��R���Q���Y �%�y3�p�>+u�l�[{�1��\�z�H�5^�[H�������c�+��J����"Z���K�<�U�Ls%��|0�Z}0�8�?�񓣅x~��cu��'/�Z����tjQ�͓�d-�.ͤ���sw�<(�uw�s�g�?����W������L�s?��������t��?�������Ń�]L��B���&��l���Cx(�����Is�� �m_nl��XB�K/�F���h=b��C�'�D�K��Y֤����zE��l۬���ʢ3g�v�̾�N|����fG�$� $�2P��{�'�_���F��n��������Q\_��I������[�h{+���%<��? �/=����M� #I2�p�B�ɼ<O�ϳ�ILc�(���	>���׈\_h���|R���@*��3���;�÷#����jGC��g��K�MdR������6X^�X4��,�ϩ\�{�f�@�I�!,�^>߼�UJ���w�'��F���Q(�)�W拒׊��n�qzy*�۴������K>��m#h� �r�-?�7���xn>~��^��<�t\<���J̷[1=�a����gce��1��|6.��7�.��Ճ�٫xR�'ʑr��l���«��v.�j�nk
�jf!�i�D`ؖ��:f74i�M����*G�Qi�x�	�9	Y!*,9z��9��k�X�ZD%RV������m�?e��F :�xƭ���˧��6�e�}�[�^��L�T���EQ���5Pw�P$�G�8��T��
�
(��h �5 �>�!����<$^�/��I��c/�J1��)���4K�ef��RA�L�5/�Ï����v|S/3���k�.xq��9e�<+r�@d����~�{��3�M��d�
�D*a:jˁ�a��
tG��9 q@�ķP�ʲ�fe9��!�P2�q�O��Z\�ލ�m�sb�sB�¹�Qv���������j��꛱y�Z<��J�����}1N�����]�mz<���AC��!� ;_��}"��3�.B�X�X|,:��c�p::}_�Ȋ�_�<�*E�zs�=c���w�c� ��ast���a��3QY|$���pР���lB~;����}��Pk�׈m��ą�~4o������'�Sv������w�b�!�V�zVۍ�#<�
)�Ay�
dL0�uG�n����"(hx�y�TZ*�δ�O�3�齲nT��?��h�H��ސJ�T����Qk��\=�u�2+����r
S��$p��Ql�����O��v*�o���=�5�Q0?/�;R���K�N,d3��H�g���mG̤�%�nJh����6}*b�8n\��~�a
Xx�����r���C��V��L<�6���,E�t�G��=��Q*��!:�ǎ �و��f����F,�OG��2r��.^�����X��4P�$UD-���R�]={j*z<�{M<$R��rZ�V�k�M Xk���l�X��O����
�A!�q�Q�C�18�E!H>,��Ñ��L����{}w�g#�.sih�����#!s˦}J����f�a�#���wp�N�&�j6=2�N�s{�<(q����_i�%$P�����rX6OS�f��s*��M���y$B�W�h%}v	�g���-IU�Wh��|Ӊ�_��R�O�.Lf)���i ��7���g�)��2��V�ݔ���2�m��p$b̓��mbM#�t˄�nz9��� F\G�!�xấ5�dB�%�&a�gޗ*�o! T<O��i�7�alc����w -�������p�l��Ȟ�>�(�\���y-�����x��wa�i'n޺�b�Ɋ9����n!��!������0)0��{H���iW�,1�]��:��q�U���ﮜ�
��>,�8� �A�����r;�Qc1gy�jm���p��z�y *�ʭ��QѨ��G�����Ug�2�������~܉��6�g��^��(�k��8X�
�����E�J�*�
��!�J�2,��Jy�m�{���S�l\��߉(Ll��+����Z��y\���$ܤGK�2��Μ���|�]W�t�q'��(â�|~�J#�����`;��t9��r9[��\��2-�s҇|@>ӓ.��~����+�>�e�<+ݗ��NE��LO�d����.tp��.0�WΒX^&���Nco�Qo�'�7�{��V������[���?�V���oū�����������(������;��v41Ʀ\SP�k� �����s����7��
�A=hf؄����s��F'�kK�-)�Iw�nߊ�֕��+Q;�F�Q뙂��h7��}�Z?tJ�Ҭ�'�]T�����$���/����X��쩀�iiL+�%|į`��!�cO�2x�ٻAV�s �#J�X�K��K�F�W�$�!���p���$
%^��u�K�j,����бJ��I'1�a��X��RvD���'��6_'$�N�����a�!�Y3)����HS����7�"\��\g�p�Q>�Pp� �ؠ��t���&���Q����28G�¶h���_�Ae�\\U���0V�����c�}���'`?��Q8[��N\��C,��ݸ����ۍkW�@ �x�����g?��۫c�Q�@K�\NnD���ôV��r�,���j�Ew.�{�T[����Z	6 ?- �ߎ\���u\Uv4~�4B̣E @3������tX�B��x��|��L�ϒJc�z;� �JܿǼu����F����E���yUzQ;܉��ZLlD����	W,>�K\���� (���@Z���B;k]S�����D�����g�?�'~mc.�C��ӧb"o��0/IxfN'��W�gfSw~[4p����T�BW BQ��|�/�P�u&�%�����N�*ЈG6�ˏ�ҫA�ɧ(��3��J��l�|�Y�ď�g�ֆ|�<�
=�x��p<y&��㰺�xԮ�'�YڞL��?u�YO��������?���������������_��_�j����o���O%����7⏾�z���^���������f���G9bl�9KY��N�G�϶�a�Ч�+��t{vw��׭�>���0����i�u�\�#��C��atv֢{�n|���br�	���j�~�S� ����D�w�G���[��]�O<G1Qg�r�t�^����XR
i�7Xlc���YԷ�3��O�<�5�ex�9D�*�zh���%������8'���^p� ����̅?aʁ.�6�O�}�[�$�oڭ�sPiS9d,i�x�y!ߥ�A�v��}Pң
 ����Yp�<�y�r��{e#2z����Ϛ���tR
_J^�-^�����}���'qj�p$�)�YA�f#(\\Z�a�I�,q�GX7#,����l�yRD�з�R�I~2*�
����@;׆�r�_ߎ�o��������x����g�����x����sq�����~&}��hNc݃���i�dK������"W�J 6e��;�8��"xADi�H��y���rC7��D��T>4Dz��R���[G��9������'��^*'�
Qai�Wȳ6I����\W�`�s�]���OC�[ܸY\��r;܎��V4b��sތ+��O����S1yj1�Q�|*d����ϳ��9���w��A��F�y$�����Ln[����%�����G�<x&�z�_�2�Y �a�|���^F%��{e8q
Ã��~ �+��O*
�g6�<��|�߻RF*a&i+��B�$$�iٚ�\x`:X����*��0�$�x��'��8��]��m�A#?��S�)�1��62=��UE`�����������\~���q�������o���V|x�0^��������R櫅ڃ���c� A#e[����}$�ⓊH� |'�vi�=���:�ա�*3;�\��UܲĮ��X!�:q|���F��M��B��.�k920�1`�\;ǫ^�B�L����!��F���KO�����1F��XF��c�8���S��"�G��Fp�!-z౛lB�� �a�*&���8H�d����&�I i���"9i�`�����/=��P��4c˓�V3Sbg0�����߸dif|�T
�)>_1ȳ����Y�O+�ɂK3�8y"	�G{�.�Kz"���U֚
j�L8�W�Tբ����K2Hb�K �~6�#������" ��gȓԻ�ӵ�Z�*�]��Ue��3�E����n'�7���:V��K��]�����u�bw{+�W7�ڭ����5X�������Ϧp����i	�_q�]��ɤZ�
 P��ܘ˅�F5���(-��]�u��dow��߸n�u�ϼT�0�Ae��Z!�a/zU�< �*�Rqw�m�ch�w�8�n=����9���4P�<�vHX<�ۋ��V�v��J��hQV��Ř�p*�K3�
v�|�)NTضI)���p���툳�NR�Ց�LJ-J|��&�xH�8�g����m_L�l��<Txj�$� ��ܭ���X�����[����$���=���>LZԁG���!�r���밑#�1#ξ�洰�d9��\� x��|�n�K��2܆Fw	�&�+4���=.9�P˚�9 ��Ɇ�[���<s����KmI;��,T�(����t��{�m��S��O~���O�T��K_�;����~�����K����g]�!}Ãu��Dw������Á�e@Pc���֣>]�Hݾt2��0�̛{��%��o��:��ژ��9�����≟>���\9d���1ddW�+л����BS+�����|����+�~G�#���^c�+�	���-<91^�چ�TH���zH�S�*dAp҃M"� ���x��N���Dd�=Ȯ��R'^�Ү���C���p���֩d~~Hy�"E�S�8�<�!9s��,[�ʣ�N�{e�|�4L����9���i
�^ߦ�3.���3�M*���1���I�eh;*P�sn�Yf2	��W@�z��
AU[H�	ۗ��U ���^& 'w�)��A�i�6E���T��zv��I�5hLp����ѨK��Yy�=&��a��b�o!P�m�ތ��n�l�A�t!�f�� <�n=v�#n�Z��;w��}��!B�m�q~�dР����ho;�����pE��G�ʲ���ڏ!��q8�n�xt����u��ݍ!
0��u��I�=��1���'Ǚ4գm��G�-���T��C�����=��&�[p�B�
�G�GG�١l`�}؇~��s/��1�}]�2И�����9����8@ n��1�NK2���1 �5�B��DN"���	����d,h�D���\�E�ż��O�	N �@�K�3�7�������P�7J���ұ��È*��c�W�Qw�@ޗ���7�d�"T�� �ظ�I�\��,W��sU�4?�g�Q���9�����y��㰦��P;��]VA"�a����ދ�S�)��^�F��"���)$#.'�ע/�oE?��:X�����X�u�~�/|9���/�����ǿ�o���?���r�K��W�{��V�O9�8�J�v�)� `�C�8���u�"������è�u��B�c���M�w�Ai�}ݣ��O퓴�=*1��;���������b�7�(�����8! �n����TfԱ��q]�� b=m֤�^#j���� k�����?��(�"�_���a�S궱K��Dz^)/�H[%���r5W� h��30���D�t}Yp
^��IjҬF�y�C)�wмs��9aqM�*��H��0 Q��C� �Q��KV	�I�O�Uv=���V�B����g����W>mp��縮尤���'�f#���'�Pt^u��T{2����RH�fd
���QK�MY�vL�pʡ����e�!���	��k�93:� �|�� ��5������>�Q��v+'�^�����q�֭�9�UV�Q��o���߻߼�����gx�9�ZK/�{ �=^ۈ���ߺ��[�[���w���Feg��۫Q�Z��Ɲ�޻��;Q_匒�ܽ�qgEy/����Fxe��m�nD/�pm5Wn���g'�/e��n�������;wc��ՈջQ���pb|��N����h��G���`�E\M�Y���g����X��T}?yI�]��p�`�	��������ј��镥�\YD�8����O�Ƽ��b�@,�y�x�^җ�x��TM��{�����Ǩ��* �[W2SV�G99����ȸ��X��˵���^Z���������sZ��	�u-h�%�d7A�@:��h�2k��F+) ���[�Idf��(���>+�Id<�#뼫a,��/��A<���OE���ic�����+��{�S�X����Y��ի7�7?��>�]��v�nڮ���}4�z:T�d4�=�q�{��Z��ޤݛX����������}P������ժ(�	`��n}1���n�r\ٛ���e->W����~����8v(��rO)�O)�U�t��Lmޱ{�38�^�Ӫ��<7�ϧY�w�Ɓ��7-i��>?)D}�?e��l���n�8�纈�?�p��ty�6o|��%��,�z7��SN�ݒ�4�0�F�2����e����(�O.�%��J^Kv�����'�`y�7+�4�&�	O���nVC<ʋ.�Uv.��f��̿����y),��	�R�-�����@������]tQk	
���1ʂt�2-�M�s^"�Mʥ� \�5��s+���^�g>�����,X�F����n��`�s�~Od��h�꽽x�������;j4*13W�����j���R��gsY�������8v`�2rTLo�ǥd��b�.��ڎ¸�Gdh�i&�b���3�wv�����\�J�P���l���A�"6:1�Ӌ�A/���xE�xN[;(V��v4�X�&vw�����n��(s��R;Q�S�o�\�5P���F�Ӎ	����v#&O����SQE��Ӡ����k�q���Bֆ0��ܡ��Եs�)��1��4Sg�sb��a�·�D���K���A��ը��
��P�B�<9!>��w��,#�`,�J1=a��[�GA�"H�X^�2d
	� a�痞�ω��i�s��GpȼE�R*�qD�kȞ�,�|�ye�^��a	ࡎ�_��!M���Pe`6�pf�8�DMCл�r�"�iL5U@
H�B��3fP�pΘp��\��F>U�hԡ�[�����ϕ�[n�Ё>����������r��l��|�����W�0}�%��F���zns���;x��r<��.�����6�[x�G�m�)�{xJ�H:w:m�qu:F-��i�����!�b�h�JP1�i4��¦�����+����q�:n�����9K[ⅶl��Ƶ$)2�t��Mxi+��H�2�EA^hJ|�n�\rG�l���0�J����_��JJ/��æ%�
ٔUF�A�w��qSO/^�Y����?5��Q�!��F�R�p_Jn��4*����%
�`=���{{O�X�{s���
�fT�g,���u������qΒ��L�)��r�)�Tz~��SA�����Aa���(�KF����%ؔ�(��.����������;���_�|,�>�¹r{;�/�#ۆq�����u1z�rj1Ν^��Ks�������Z�� �=$�vp�-/���6MQ�����{����{����syF n~'��Սwr6.�h��& �	�4|G1U<,�P� ��
�]"a�*�� ��{Ѥn�ഁ�@��\������XV��~<�ȧn�X�Ei,Ee�ʻ�=�}�h�H]�X��qp/��f4��­O6bzi6������!��K���(��&�c�`=��}��]��1A"=��x�� 	9[��0�)��+��ۅA>�,m����͕�s"p�0��~����3���`+���ҷ���{ҨDsf=d��G�c��V`�D]��@������Y6<�Z�kH2�'��
hP%TճQ� j�T6�@�ד�-,�Je��M�Y��BH�v�Ǉq����ٟ�7�z3>��j���7���69��{ ~�_�G}��A�b̈��������[x�ݎ��&��}<��oq}=��kQ��FT|�G��Z�u�h���u��eU��ތ���A��D���Υ�eg;�E��B�m�g�����v����ޤ�ك���y0t��Ic�v�����>�`�{7�c��� ����fi[`!�!|X�a�{���Q�z��{:�������ش��Cł|�Er�g��Y��I��Y(���!�,�;�
dJ,~��M�*�o��6��,�l]i},�������
�I;<�ہ��K2-��2����IK�A�S9^`3��zE���(���WE��Yy�i������z���2Y^y�8�W0K�d Q�BL�'�$�n|?�5)�� 3�R3Cѿ���T��|;~��_����g��=A*(N'
_�0P�̲�������<�w�}/��?��������k�7��~�7�o��ߍ������_����˯�^��T3&�+�OC���#�N8�rٖ�&�?��{?����k�XW=�.��u�QB��P������u9َQ�@P0��dZR
_����H-��|�,B�I9#�����H��:�l��{󷣉�3u�ga.���>D�� ��CP����x�X�C�
o��էph�s=���ә�!0��~Hwej������.����T��w&��ٍ1���97�_&�J�`�g��	j�'b��ݹ�q�|k(�eM��ľ~�`��)��*p�G*���B>K!�p'�����.��W�t���MoHeQ�[(�p�A�UI�zzz�8~c��;(c�e�#�XOꏢ�5��*y7)�]�H��e�V�(�߬Jg��0�����a�8��>F�C������.��S��0�����[م����Gn�s�J�UW�Pn�A�܎эU��5��!�VT�PR��x�x�x��]%�����oǔ.䦞�����~'j!?&��%=��OL�"���]�������>�"�B��DAq�/��zM���B���F��a�\��jpء��K^�eHu��'��Z������5�J�lD�A� :�P��q����S�>�2h��� ��  ��IDAT�;")7m?K�',!o��n�'e~�;��T�#o=�F{6��R&��4в���2Ձ�҉@���8�|aF�"��=�d|��>�x��A(TR���qJ �s����c�<<������ό4����_��{k��_���L*��!2v���>yw����������t�dn/ʓ<d��~��!ֆ���������V�x�b`�Nn��yL���Y����y�f�ݽo��Q���G��6{/��ڏ�.njs:VV��C?�?�D\��R4&]m��;G鎣�:�����6�}kv>���TU��*^Du
��Fq����Qh5�k��4�
S�����4
g�eP1��i����^�f�2����yDy��6��t��u>��ʭ���2���,�2k�
��lY�x�3�2u�G����ʰ�=<�lp��9��鍍�ov�� �Y���c��٘X^$�Z��� �a���q�./�0�-��I�RO(/--�5dN�����f��_�X^�/='��m����8޹� @�ډFk��0x)/9�Ԟ(V�[\)�z�I^�4�k��M�^UzNcZM�:!8�H�2fVL��&=kk�T**'�����[�u2.�Q^��#������ y�٫��GN4F'�/��@�G9�V�]��Y��Mx�ҽ��2�K+��c��T<p��8�\
��z3�[��|�9�kyy%Z����� ??\!��]�᱄���eIdP-��ˠ-7d��OIzq��������(=*����s��C��<��Ŋ.f��5���ଊ-e��s,����8�7����/Q5����(�k(���x��R�|�zV��6g��9�l��������TlE}�ӓØ[Z�ɹ�1�h�.�����?��l(�����f�ez��)qe@��e	�v��4�̒�\�!<<��v��h��;d4���2̜�I@�5nr^
(G��ZE /
�L��iL/<�I��D�y���M�~3v�����:�w<8��J����?yܖ���3�)�
����~�W����^l�
7����^7��۸Իq�����%�z�a�!�N]�¬�c�d%?�/"���ߍ7>x'>ƭ������j�v%�El
 g"f� l?�����t<���3�~���d\<���cuc7f�q��\n�u��t_��Xo�o܌�;��g�܈�^�F��֕y,¹�[�2�]$�:��OJ)�����
���q�����7�s�hx�[�Zg��N$=��r���-����׳�֥\-�݄��(�Y�_����1y��B���^�����z����Z���M<�N4QP�Y<�s��F��W`t<�}t�~�>��УT<0n��C��x��؎c<#��Oo�۳2Ѵ|D�Jq�'��A�]� �]�˕-Z��设{�ތ&����Ӿ;�S����6��9�j�_K:s���K�D;8�N�U<�0r�cv�h����]P$��6g��K%��u�\��l�"�=��ZD���w����w
���lgNE�6N(�8Ѵ)��L�~�rQ�*� '���? ;ox�|��I(�~������B<���x�������'(���$���/??�s_��>���� }���Q�ݿ�;�ﾒ;s>����O�T���~;=�Q�H�b�Ҹ�"����j��)��%����u�J*-��g���s������Jm2�]>/��h�����<u��ﮫ��b�ɛ���R�#�=5?�W>�|,���b�n�/�3��1���1����I|�����8Ӎ|����g%�O����q�����P��Q�W<�����d>X~(:�y�Y�J{T������Ӑ 7'���|>�N�-S��]�ɧ�vS~
�Tz4é(����¼,����W���*8��Gc���<�W;�o� \�����
�ϥ�TV6��r��H_z:NV����=<�#e�=$+p���I%��qs�t�ܸ�2�W0p;�����S�q��ro0#2TƓܝ�k_��׿�����'o^��_�²H�hGDčm����*��#7�S��dK��u�)P�ʖbz����������w�����@��*އ�P��Ξ���Z�駧&⧿�H��_�Z��_���җ�?�g�L����b|���ŗ>�d|�����'�x0��l,.�1� �N�Dބ�n���n
(6��3�^X�����cE���6�x#���5^nWy�Y/��ϸ�x��k�#|7���C�ɠ>���١w0KLN�gE�I�ʵ��	o���T%ވ��ߧ���1 �A��wY�I9�q���|D{���1��$C��Voߍ���h����P����1u�tTV�C��y傞��FZ��Y�-�y�&?`t��폱�nA�Y�,��sW�u'�rN-ßYi��mhn�|��Ԥ�\
	�T?FIn#w_��V-��KX�K�;�2�:92�L���fy�����O�c��oE�OGU�\�X~%��+X����)]���Q��ʘɔ�F�Ӎ��Z�i���*-�!Rcj&��#�d2�/hd�U| �zM@%_j���^�5��./��D٣M?�oO+N��ʕ�߹r+b�F�d<����瞋�Y<z���xna�\\~��X]ی�7n䢠�z<��x-*.Y�}X�@=��`<�?O=�|���2�oO~
`��c�#�̧�+��=p�MB{{�c��G�����V�$.J�@����؈�u@!V�m{��Zʯ���8wy%^x�|<tzg12NA��{qk}#j��x]��_��ˏ�/<{1�=2[�1��P��UЅ���3Q=7��TTd���[m좧�M��|U�ū���A#WHqe��4�M1�<�l���yTd:��ƕ�g#�+�B�S��>�B����U>��>F�;��z�r�vl���%��<�}���`��T�	���Γ��k,�$(�+�CC��B��(;�@V�(���#��B���g�C��s���*^q��({Zx �(S��D%�x��3�����no��|paFfM���/�@����p"��ƿ��/"�܀���@y(.�i@�uOv�t���ۿ�;�+��߉kW����e�o"�!Z?ȶ�zCu��LƟ��񵯼�<�P�?��e7�ӵ���p��Ԕ�|�:qt���0l9O�=X�7?\���<݊�4B���F+]�>��R�5�<� ����D���N�1�,F0�\O�`M���s�,0nZ?���U���|��=�~���GY�7/�u��+l(OF��)�!8���;�>�+ې�]�h��x�Xo�E��V4P�v�M�[x���A�/�!Lx ����X�dj��%K�r����v���A�����}<<�ƌ~0Q;�n�6��B�"QZѣT���#�,�!�<��8>���3+@���{L����XXZ��r�#�r����	-�0�^��I*�!^�p�����^4+��`s���MQ�����X�x��S�$s�m���h�4��nь�(���"�1�wqh�,�L�+O��޼�b���E�Pπ'�ॣ��0 ba��������J�}�vT�n��^|*~��Ǹ|�\���;���O�`4ǅ�K�̳�O=��Y��8s�x��1:B	'C#���3?�����������g^z)���PL/LFs�G�C�9mSAID�V�zg��ęӳ1��t��
�l,]h����X:���P�gxw��߷�h��ˍX�8+�fc��r���//ƣO^�GOOƫ/;޻�x��7����6c�]�gx����8Ё���x♸�٧c�`'n��p�!�F#<Q����^�]���v�GGpCs���U�ѷ@��\=�yp]�ʗ\�1�|i��6��1>|'ݥ7�-����B�^�k��2���\�{� ��v�?&��Fs�p-G���<45�$9V>�g�BHX��r�8����F%�2��k��nw7����TzT���L���*��0�G>Me�I��f�f�0��n7hY|d>�� �����n�����~�[[���a��DZ���vA��/e0a����z���E���?� Mh�]
�8w�/���k���V���|��Tb��g��0jYa*�*l�cY���t����'�/��և���l���Zt`�w���XT;�����q����ݵ�X:u��B��3��hk��W��bEy(n(��� Ԛ@*(��
��A��*
&���q�|�t��3��јrN���stZ����Ky��]B�˳�X�����i��6��ǷP<0qs�(7=���t�/-G��".�D�I30g�s���Q����p�Bl�.��߈�ᵨ�R�V4�/�-M���������9r�8(��rԘrޑ�T� !�:9sgû\��.�Q��k�����9J��1�LDYM�<�O�y�P���k0��������h�L��,`�˪�0�"pRPd��6�U+}�~R�z�,�Š��]������RQ�ҶZ�BI�� ?S!�݂'��4:S�����խ�C����,��뷢��I������K_�����(��*Z^Z��9�u��[7��Dc
%>��ɹx�Տ�N��C}%�W�����~>���+����xn���F@=��~�]}�6iG����7<���=�h��G����g�y&>�/�O|�3��O<�}��x�sO��/=Lx��@|���g_z4�}�x�3O�����^����x!N-�cO����ym�V;Ȳj<�¥���?��X��O-���|<q�Ÿ{�v����})��"��c�w?��\a�..���=<�0w������V��V����Eu�����B�v�L�)�J��CZ�y|J�>J��QH/�,m�$3���~t����T4���Z| �S�h!w\U>S2��<�O�$UGfkv�v�u9����$}�~&��EФI<��M�<%���V.K��g�F,
M�'=�n7�N���Y#�ǔ���>s��������W�ދ��G�\O���G ��`��Q��7�_���ᭌ��P�wbbz+����ߊ��n�f'a*\��kq��G�_�׾�jL��	�&�����+XzY�]jO��'��C��=9���U�p;6�������z�ݺ7n܌[wn�͛�s��?�7n�a1L���G����p{��|;?؏\��-��:l�lHJ�.֓ �jI��r��RQ��F��X6��Qb���iĲg���bE�DL�H�g��Kp\��TJ<�T��	���ґQ����V�n�GOv�����A�3Ѿ���Q<�ܮ;#	@��j�O���(�j.��c�T�2��ۘ�Ay_�9��E���(V��E�&J��!��]�r���g���U����)h�F��⠧w�H��A�+�璿�����CT$0(NG�'-5�r-.���5u坏�\km<"f�|l��9\�ϵ�dbz ��b�P?W�se�b�P+� q�@xK�țҺ*Pў�S)�Q=��/�`�w��!��91w7���313ӈ;\ݻ�P�c��,��a����,��s��Vܼ�Q��?����?�>^f'�6��^��޺B�*��D�9�D��_�\|�)<MʷO�;f��Zln܉G.]���/������?�`���})��_�����x�y��s���x2�|��x����G�gx0�}�r<���x�����3���3��3��}����x���|(�t)�Oe����x챇����O��Ǔ��B1�Z��T�w�?	���������Kx<�D�|�3���Im� �H�.�Q�)��{���:�p�8�Ɣ�� !x��\}z؎��#i3�KDiGS�A��H>89w�\���@Sgc4�4���
���ݸ�Q�W�R��?��<���Jw�_s�K��b�d�;9\y"����o�q��5w�ř�'�-������T>
्r�Kd艬�y	,�(�ڿ���o�܊�}�.�Vf�;%#9�2���F?. ̆��8ڽW>�(��b~z.~����{��{�r���$�b#��o�Z|����ɷ`��X9:��b�:e$EyV������)�?;�#Rd��?z7n^��7o����qo}5��و�܊�?�(^y�����ފ��ݸ���
�������V�{���C#O4q=A�M<���IZ\g �r4	��Q�l6@Ґ6{���}/�e~�,q<'�}H�r}wB�c�杄O>4D�ټ�~��3�Q�)u;���\P����q�4݈��\La��O/D�!�zjR'�۵�,A���`DB��M"����������NeW��Ѯ
3�����5&��MUɋrT�C-1"ro�z��G��[�g��Xg��C �<'����ħH�ol9�� �� +^�K"��#Y`�����ີ�8tD1�IԬ��8K�e�R���+���b81Gi� �#�l#���%	'��Bx�m�/)�0WqHϫm��ӗ��s�����y0w7�ts˳1=���7ߍ{[;q�ڭ��ߎ7�|76?� >~�����ߌo}��߈�>���c��鋏�{&��[��R(��}$~�^������0�����wb~~6~�g~:~�g�/>�T<����?�l<���q�܅XY:�9�unv��٩���S�E	����ٖ��܊b�efj:f�=Oe��ť�"�:��$m�S/>����'���S�����NL5�1GY..�7���}����^��D�Qe!��R��tʯ� �5x߇l��F�#��Pr׫�,s[z�ŋ7Ox�ǉз����c��[�S������z��C�yP�)Zf2:hz��s�ge�4�B�<2��(^�P�n�+��M�Q��u,�yg��%?aOL�ߥB׳�yFER!e\KT&�ǹO��>�J����3s3�_Ҥr-ٕC�/��&�o|���x� ��k�P>]*	�x1E��5XV�{4�f?>ڸg��
��G����݌o�ɷPD�ᶪK��q��Z������_�5���0��ت.F��2�}U�# )_�e���0����o���Fܦ��x:;X~{�f��t��n|r}3�~�N���'xAwcw�%�۱_���7Wk�Qrj��9�׏cv/�/?\l����Y'���>T��8|�<�r"(��$YҘ>���&��,�>��ÿV����=�]<7_���;�<$���o\�0:��|�j|f@�D��*�nA���ڋ
J�����^�t���tK��b�Q��Q�d?�����]��~S��^�`i$��=���Z�AE�"pi��!��f7�Onn� Y'��L,��O��h���d�
�#�T�Q���`�u� �.�=�Wf�J� ��C�l��ޥ�L�"�hb.�X�G�^Ov:$,YW����<I'J���n�J��
t ��x�*��*,��Q���叅O1s��5��)q .�6����^lB㕝�T>ⶽ8�x��8���o������ʝ���q�V��ɭx�k��F.~��1n�693?�d����>��� 	?a��ʟ�l<t�tzR5����Zܻ����|�� �jV���p*��v��x/� ��'��}ȟOKہ�l�77���o�B�D��ý���_N�yO�Rkc���
�9�أ8<��������?�%���||��Np����^T
&ȵ݄MC�n]گ)�����a%,�x���Ǔ?��6�"+nN�g�M�G��TYȖ��F5hZR�����	�����3/��k����������U�[���.���H>#C�O2�^şu��q��:��iA�MZ���=@�y>S��N'Gr��̓#�'@�U>_��׿�&��o�q=:���M*#���:��������Ek=�����~�oǫ�f\:5K+g�X{��o�w���b��N,���϶�9����~�� �t�˥�Z� 7t$�V%^ʇ7���7?�����k'����KwT��A�>V�.2�i��Cd�(g�w@���U2�A4�t���{�1��G����Y���^�p�;{q����~�{�{�ϵ� ��K�8a�ᤤ:��|�#�3�zDy�Y!N���;<ߍ �
�T����ky�Ý݌c�|o>�4$_�n�׆�F��X��͘\�
���sq��y a���D��ų\�&���Ѓ˶�@�qPP(�z(aPQ�V`#�(�	'���4��N�\�D���d���|��Σ�}� �-8�wht��QC(�B�+{g�^�*��҃��{�hԄd�&�Z�̜�����l�d���T0�4y��R�!��@��|�%����s~�JA!����BL��}�s��T:��e��g�D';��Q�����F�V�����l�Z����alo݈��"��w]�Ɖ�sQk�ą��G5���\|�s���v���p~R3f/�g>�H��V��z�Gqo�N|��qk��D\8s���x1�rP	� �d�l���XPe��S�[�sSRpϵ���J���N�M'k�������z-�\�2?G��8>�CNm��ݵ��ފwo�o��?"'�:ʧ:��Y���<h�~ı��oN.�d�L�c���&�[W�+Z�u�K}H)���4'��������r�y��l���/�K\��T����#���K�v���(/�3���'=.�>_���Yq ��6�db�9��ty�Q��Ŕ=)x�M���v����59�E�e������wBW����< �����o|����ۯ݊�}=
�rD/�,m8E��Zi���+��z3>y����ko����0�]_�~���?qp�ߏ;wn���T,�����V��<jƆ���'`�P�
�S��/��ٕy�~��Ļ�܋�~t��[�v~m���9�Río� m�%���Q��*�B�u�V�m�;h)נڅ�]Nȕ�9��˳}��U�}ǹ���΄����_(�����R!�N�<�`ԝ���œ�����F�y�
5�RVAb�|G���޲q���Uw�#��G�ƭ��~�P����D-=���x�g��;��D1�M��(=s�O��lj�����,<s���J|ڋ��B�%<�����
]������kOfR�e������<�]= �d�ӹi�k�e�ʞY+�r��
�d��@ϩ����0o���܈�s>&��9�t�s��;NVsp���!��s��`�X���^a�Bϐ���.'ĵ^���L���:�G��v� /X��[�K���}�p?��g�>�h<����s�ǋ/�d<��K���Oė~�x��g1N�Z�ٓ�r�L�]ߏ�OTU���x�'��y�����������;]����������r��.�igk#���"�r�C�AU7)��8��Od
��]6M>.md:��^o;��y�\������J��p"���s����Nܽ}'>���`��`���o��Bn˔5qz1b~���WidP.�!d�/��¡�����z\�T@�������lc��95� ��^�hY�y���t���s�J\`�p�+�Kߜ5��³���-Kڤ�,���xٽp�'�x��J�lr�\�%l$I�]�)��1��b
ն0��@�z�:�v�] �+���':x��37�,+��0��;�;��?�����j��`��0�&��A3�Ks�X��ޝ�~�f���1�?w*bz2�ٽ���4+�����
:�i�O�w�eM�	5I��@K�iG(��]Xj�\�8ZXE�Վm»S����$J�9������Ԭ�(��������^�`1�Z��.���\�2�=��DFG�V��<3n��=�h�9��y_5�
P�^�&���Ƚr�v��`�T�kw�����2�� Z�p2.J��*��g�Ui��uaӔm����BL�tj���C����t���k<K����d+�/y��d��1N��.p��h��Ћ
"��l��H㘯?ҦB���3�r��ͭ�����}��n���~�Ǵd$�C2�A�)�/
L�{n�I��ģR�
��ȱU��r�-{2B'�ܼċu2?��}~���H���݃��o��SK~^s���Q�=��C.���t�%���j�}�~�\$s�eS����;ݷ]<�=�h����_���~<>��g�_x1����'����g��whee1�~���������-h�S���cW�w߉?��w��F�����i��S�|u�[�xH��J}�e����Q���E0�ؽ��E�Uyn�&�	�G�W��6:f{�?�ַbs��Ξ�6�feЏ=<�u��ͭ�ț�_#~����
�*<�9�.j�5mB#�"��]������Ю�g'�IRҒ�M���	2�y��Jr4���p�o����Gy�lk�\�t%���|����*�\���<O���t>/���#�I�%{d^cp��X����'>ͫ�N<��C�v�w��, ˎ���ti����Sm:ާ�q�W0΁��N�k��q�/Qz8�p<�XN|�삊o߸�[�؝<=�KODo���Ո������]��[�)�8��6֌���`GZ+�%�������h��杻�������l�-/EjX�"}#-K��̼�7��,��b�i�7G6͜�҄I&,�����J�u���Z��n4k���kԸ�y
TpS'R
V�K�U��
ξ��K�K��L��3�-�\�<�A)��m��@�H����R�CH
�B!�ыK�;�
�/�65�K�4�-G�ҙ�b�����/��hy��6|�(�b���ZI�F�k�QO���	�����&�� |)lɤXO���
�-� �9��}=��C�#�rɼ�	�4��,;��x�w"�?� �M��s§C=	'މ�S�p���n=�Ws8���,�.$��a\����wz|�?�<���-Ft	k���
I�W?���<S������ /��v�x�E�ي��L��W�L<z�l<��{a������t�8�l��a��p�\;ΟZ�����~}5�AG^T |�w���މW߻Wno�-��i�@I����N�|
����T%%�3����yV�<8�ⳮ-p=?݌y���^�bԮ��J��Q�n��:�?:J~ҵ�.�2T>U��k� �=�2�m:�I��k��/ʃ��^�6�Z� Nτ��|��$�7>1m�|�+.�!�g vC.�D(�Y�́Δ;�+*TVx��GH#HR��}�KPRߤ�A
�IYc:R��9���?�0i&7߼�<qG>�0>��u��d�q�K&^�̓�K4�w�o|���x��n���X<X"'��eDQ�K
��=�wpw��1l�	p9v�&csw[�Q�Zj���l\�܏����Q+n�W����9I����2�U�wb�z(����G0�}<�^=�Q^{�
g��h�"�{{�q�v'>�u�V��32ܤ�� ��d3��AW�jmҶ�Q'�"v�W 0�4�)�y�a+��U�V�c�9L��=�&���C��{� _�e�Dݕ�A>����P���x�\ǭ���9��f�[���y��"��q��OG}y.�s���tt�8�N$b���*Cy%S&'�����ϳ&�l�Ԅ<LALPh�b@�������<Hw��$&�d6��=*���������2$������&]��{~'�̔ㄠ��r�H<R3��
e�D� ���J�����a2���DQ��h	���,�k������>֞#:�B�+'Ц�q��T@בܭ��7?��4t��q��|,/O��!	Qd;qx�xH=��p� �$lon�����F���zo#޿r+����x�KQ��TL_X��=9�����A|x�n,-.Ɠ�<���酩x쑇cbʕ&�i�:�d�����u�x|����:|&�:��#��Ν[qtp��?@��t�;/��ԍ��;gN��{xc�{�+v��'Ũ���;��t��x��bn���?qL��S61�|&�f����T�	g�$o��J��bl���44�͗�2)Ś�(ӕ�J|d�c�%=����yW��Bg��$��/喌�����]�_���$<��8朹�0����8z-��Ʊ>y?>[/�90먛�=�=�9���/�	*�n.��Ν����|��h����H�\l��[g�pxX�^�<@h WKn.��k���/��wo��[���ۙ��C4'��`Ԧ� l0�i��~�ֳ����(��N5:�::�\;*&�q��n\�qa�w�S�S�����i϶bji>��Q[���|;�s���L��S�몣.ZC��'�VPƭ��g'�g5��<b�g�xf*D}~��,o&&�W��<�ϮB>�G�+����w�"%���ܱ��`>Iӷ�/�A��)�&��ʐj�c4Fd{�<I�R�g�	�h!�Lk@)���>d�dҌ�HAo"�Z���D�0�Sa�e��Qј��B�&7O�6�L�3�ˬ���d���aYE��g�0ȉ�@����{�ɻ
˱>),�{�(9������g��3�3���$S���sqK`o/j�ݤ���I��\#���E�I���g���m��|4�чٯ]�$Vo]��{wcw/Gu	ۤ����w7����x����w�ś�7�*<�ׅ�F�F��ť��g��3�d�Ϯă���T�n_r���Gs��<1{�[�逖���G< ?���q�.%��ы�W���<�Z.�u�9���fl�ƹ�1;3���L���?��'} k����q{�|�1�r�iL�h"&P2����^���'}G��F	�'��$���_��I����_i����x�u��)MWβa��>�̧tXd`1�#|?:Lm^%[���k�N����Q���M"��GG��w^�_en%˂���(�
��i��^�|�%a��c�X&����v9��<�D�P�Q���@fn��-���n�6T<�`�\IVk?��6���|�w7�c�s��k iw�����qh�n�c�	C��x<?�b<�	�"����Dta�k�x����F'6v�ρ�4��`xSx�x	�x�g��yf1j�棺<�Q�=B���\Q�� ��!��g��3�^���NM��˘��5p�}o��9Fa�h|?"�Լ�(��?�~���g���������g�8�Q�a@����^�؎�u�Rv�t����e{&��~zi�I�����I,^�Ti��(������\�֮?����3�������9�g�/�A9d�(�h�+_%���||w�6	0�+��$��g�ʚY���U���N���U�����I��$�T�����R�ҝ'p���K%e�L���7��t)|��~��VT�ߋ��k�߉��Z4G�4��м��b�%�S
�9��9�kۃ����������n��V��wsg+v:���k;q����zk3>��w��q 4j�@���h�P'^�uB�
�̜�ig��Ġ����s�}�������#��Y�3Ў��T+�f~/>�tS�<�,���>2e7��삟D19e��-���mE�	״��F�����8Ƹ���bb����o�<�[���",�K=�A.����s'��m�{Jzehn�-�H�g
s�h.�u�34u:�I\ܴLgj1MJ�'���g!��o�vrO Q�rx��W�	��2I�t���|��'�.śh|-nơ�>R�5[�C��S��$��i3ss�̷��i�dC��:_���H/�q��Z]�nŃgV�Ts"�P6�8�{U,�
��i���q7n�A0��ي�I�|�݈F���|m�c�@��D�6��y�	��,��\� �gW�b��8��?��Bx!&\c�g3�c
�pKn���3��_NϠ�]ȱN�C�C�qn�� �k���C�(J����:�"\8����������o0�ߧ�T���B\�G����~	5���?���a�����,k��4�xEC{���V����� �x�=�5	��o42@y��uI���d�Ч�8R�!�)�����ڙ�i����Oj���W�q\F~��Z8
c���[�	�'���LZ ��C�
��9�*�O=����>	�f�U�P
̏����?�6=�2X�JGGe k��DBX����vt׿��oG���]�j����F5�_hk�� ��>Y3�0����c�u1�l#n�ݍ���q��^�^�`�uc}k?z��1ϣ�ZN���hM�x�+:�N��z~<>��
��]��:���C�/�ɺr\�^y�?x�t'�t`"�����rދk!*�Z���๛�Z���V��F-��~F�ؖ�-dL�,t��T;�N��e2����޵hl�����h7�Di�����K�����_Z+�ͪ���((&$ϴ7H��?�Q��|	�\f�/:m�wE�Rz��A�,4ft3)��൰i ��{�sl=��.�"ݒ��k٤�CWI��G���8�{�^�#R֑�T�Y�Q���� kK����;��O�ܧ��y�D�p?����L+汆�h����g!�Y���L=��qjc^/c&��Pӱ՜���$�b%V.���ٹ�;u:�V���镘"L�^�#Y�ƹe©h�_��9��]��yǅ3Ѻt6��3�����31}?�y6�t�?p&�<�g̜�|�xgb�ҩh��[������@8Gn����1	�g>O���"k��L�(�h1q��E��Md�HS�ƈ�%}h4�!Ҫt��2���-�X,�V���#	G��ąY�����jv����y�����6��ڲ���f�'!�,��=ϋ&�8Q��7?��D+���\�-�u+����pO�&3sN,�l(7���`������ɫ≳5T�y�`D�.�OB��S�O��O��ע�
�<L���5����yf���=��@��2���o�C5���1����l=Z�w'��GY�gIF�3�k���cQ�"l�Gq����D,�TPN�.��[�ƛ��{މOnl���ǽ�Nubb�"�kq|�nT�ݎʝ{Q]݉���\^A�[�v���;���]��>��S��W��v(q���e\��)�F���	��O�&�a�I_����s�-��cꃧ<�/�\E��P�a8��m��CQwQ�wcp�1���ߌ���j��9 I��JdI܄�qQn�����<1��aY����8��ԘHCB�U�ָ.�🐸  �����v%�dW�~,?:�+�w�[z��Y���8�^�-<�����IHjWuS�D��(��h�c�R���v�a��Ŝ���{��+�,�(I��e��K6��L��������h�>�v���&���	W˼��fmx33�Z�����X"\�#����X<3�K3�X\�����;�M}�0=��l��_���U<��^��C��j��4<���-ȧ�i��!�Tf2���=*t�U�ж5�W�L
�"sh�Sیυ�2���i��Q�Ҵ��)R!Bӝ4Z
P"'��Xs4����3�6���07��$a��oL<{��I� e�ϴRr~�>��׸���٘/q�M�m,��W:S,�H8�"8 &i�S��\��R^;�Z�t�JȲ,�L�Ώ��ޖS�+
 oDs�{+L
=�JʖWy���?�}��z���%M��!�Z��]��i!�,�w֠*�,Yf�aZ��/fLFc��p�v�w�u���h/B�O�q��ўB�GAs|��� �\n)4����Zǲ�����	}0���kO����f7^�`5��֝x�����6�����)x¶9����c?睍V�B�f�>[G�ڛ��n�w���v
�(�*��Sks4�B1�Kl�8'G�Q�������Sv��邥>ģ���C�e�:dxi�;xl�X�����;۱0��A>��
{�%{���c�A�W`�z�V�R���fDg5��wc�ٌz�����y��[����^�4N��*���By�P�I�J5��#[�LZ��m<L@/�.�e>$I�}
�����g\�����DҐ
Rn�8�^��La�"�3��o�7��ۢK-3��x_x_�w�[/�z��5� �"S�dޙQ�
U��՗���$��k�;8�#;��C8�;p �nP�h"������<J���h�}K�qyy��A��]I� ����ِ#,;� ���롄�;�*,�g�;�Q������V�.'5�6�廜��� OK�`��0C2��P�I|%n�y^�I\E�{���3������k5- �LR�a(��(oñK�s�UFĵ<�0�|rM�93�d⃓pSF��,o9@ov�x��EF�X���{P�>��fl1ȃ��ZU�5��ǅ��	��	e����3��K�'��>��gv������,������8#'b��0�?�z�Ff?Qd�.y��"��k9x�*�*���c���D�-�C�Œ������n�D �&�0�����1�|(��W5W/vpnf/��3Wv0�� �Mn��n����VL�D����A�m�c�k���t4�����8��}Y<g���[�%�5z�~��r�w�bL�����[o]��w�����ִq5�8vҦz4u	��J���O��7����$~�Ib��.ǳ��f����D_ @����!�Q�Pu����j���(�[�1�P�=5\Wu^O�!�<�]DS�(�
r�1�a<wC�|4g/� ���C�)�4 n�Q4��1Y�-�փ��t[*Tj������@~9��y��*ׅV�6A��a槐,ÿ�xɋ�1�'_
MF����g�r�T(�ǧ�PD����99�4Z��W�'�Oy�{~�'��G�F&�	�̠ ^�IgĄ�>�!�6@���J�8
� qt{��a�=�e�ܸ�9%!u9tW:�����V':f�.i�]�1��c�C�x\Z��.�������}���SΎ/G8{�$�sVـ���R�[�S������\�E��H����]�Z�.�u'K#���ނ��r$P㚞�(�䊴��6������+�\R��9t���kJ� S����p�i	�E��e�m��W���fY�e m)<�����/�LǑ��>���4P������'=%���A�c�}"a��@Ǐ��2T�GQN�t�Ha��>�>���G��<���|_�*�OX�/�%w�Uz��4���S�O�q��M�R�+��W���h�S�g(g= m�m����b��t����é8��$�c�M̒5Ŭ�u-ɧ#wz�q�^����q��a�Y���A�ۯ�Ȧ�3h�n���jl5QH�׊�����?AyQq�tgJ�Ѫ���d<�ȅx�3(��������[ĺ��ʬ�GEx���FB�:����*��Io!��+�%LNNƹ�S(B8bi�Q��5ь*�a{k#�_�͝�8����z[�l���̕#��'{��z;0�M��꼱��0�vbf!��?s~%f�rTg/�q�v�g��X
N�!�&#�W	�x��P:JE��?�Nv
qq�C����>+�,\j.u�b�Ce�|5Nw����81s�o%���M��@�XJҌ�[��[Y��������_�A~r2��2�zd�6q&�.�/��i|�sc孀59��x��l�"H]������)Ty����ɴ���g��}���x�0>X���1.���on<g0�7B��ZbT��GiuQV���O8�C��T��P�$-Rp���뜁�</]Z�C�'�J�����"�`:�-�T�)�Ń��������*�{K:�Q��d\�@��E�w�J�f�J�U0n�(���G���it��������t%m�x�"�#`��	���%a\�?�#�aʼ?-[Q	����ҎK�7�m��AO��0�?��ɼɏkqc��� &|̘s�gI���C*⧢&��E��|� 9��W��G�N���JކR�O�͐B����Okr"�P��H��Nu.��]�kx�:�q�֙�d~�����q�lw�+��޵��d�8�����Mb�50�Z�T���Z���6J��v-��q�i�������ѨOD�rj)�}�R<z�w��k�~?>�v=���9���"�ZS�������y]nEˏ%���n���:JFvV;���C o�>[��qw� n�ٌ���4ʺX�3�?�-�d�zA�ņ��J�:9�Ѫƙ�V�=Պ��^$���Ř��|��#q������6�Z�R�jQ$Ҥ���3qF���n����W�O��M�S�ϳ��+����%���7�#�*���&��Pҥ�u#�w�ɡRb�Hi�_�_�-�7�&��7q$�r�a_uuWuU����}�{�A,A� �R�E{ƒl�Ȗf��%[�,k�
G8aEؖc��<I���Y9�I� 	 ���������}�����9}/(j4!�rvg�sr���/�%3O��F��$���x#j���Tb]v]O>���E�E*u�f�rP_+A���������p�\�@�ܩ%�PQ@�1�H�G��8�5)Q�O5�r<�L��3B(�9l>c園��tgO	�ڧU3O�}Y+1�ܧ��d�����n`l酓g�*۫�\�P<ׂ+~j���`�\��e^=a�f�y�<y�W�6��&�g2S	��2?\���u�ܐ��+��� SSM4׉RH�����I��&�����O�=	�皠$�:M�W�[�
�yj��
щ�by���/RVNBvZ%�h�/�k��t�!?��#����N|_���/�~M!y�"3yRap�����e;���K�S���2ʳ�no
c�T��v
���FLN�b~ٵ_M�~��"�H�u���6@�J�6���G)y2���(N}�mo�}�C�;�F'�I�� ���g=Ka3���6��-`�B�%"���65>�[W�r��ݷޏo��V�E��8�y[[�qr|��>�%�ܸ�񞴢$)�κs왦«x�Nƚ�Ȍ�tzz�h�
�]�;���ĎOL�s/��o݊�k�����PM�F2(�3��d�>����ŕ��X^j�e��o8��s:���h�W�L��)>��@�Kň��6��JƟM-4��^AA-���xi$�5#����m�露��r%i���̶=q�A �r�Ȑ̨��`����J%��v��Y���$K��^�z�����%����/���' ` 8-����X�	1u�ɸit�C�fZd0]z�B��Z�D&"=ʦ>�L�5�oA�M��!�f�E�B�h�{ \Aĳ�D^��s P��a�L��3]�+aD���M�sU��n��>��*mAf�jLս鋰��I�	N���O�Ġ�r�m��S]T,۝�S��"s�R�6�^�)��J�-����|�"�F|�1ϖ�ŖiD#��۶d��_y�j��W|e�
�/�1�$��s�O��宔_"#u�2�F ��9�
���#a��HcZ��+���ɟ0���
����(!%��W|B���A�*���9�����<.�_vt~>�G D�S�4��9e��`NX��@a�T�gw9���>~�=���,�* �v���8oMƈx]��H��7�c_��- ��P�����plө�>	����У����h=ݿ����љ���[��tg9cm�}�������o���F��#Ev�(>f��2e�/|��y�O����=�Ȟ����Gq�u7��ߌ�o����\��O���R�]Z�g�6��x�tb���x��۱s|FY*
f&��S�~��>J�I�4�{XV#,�Q�P��S'��ߟ��TR��f���F���2M_��V�k��/		o�*W�Oz�����~˘�&q� �xY^��q*�)���>g�W.�0�Bs!5l�]j�x�)�m��{	s	�>Nز1�T"����U�MBp�Y��Kum��/~��7��Ͼv/N6�
r�	@A3r�s�. �}��C��2r���U��:�O�R��T���	D;!2©$��3�k9��Y�yE���²���4?M�X�e�+�,�R3�����'�hB׬7"�J�E�0\��_iSv�W��g6�IMc�%��W�N	�6��'��� ���S=�d�,��ެG܋�B���g˱~J��M0+�8����7:Q�ĕ�
�>�8�,����������L#Ji<eLf�$�:�)��rz�~�}x۟�����oE?6!��HT����+�a����*.��'-an��g>��@����g9��'�^l�0���|Mŭ���O^ilV��3�דּJ�;���G��x�\�*�A���D��N����s��ZNИ���i,L�i3��a8�33%n����Ϧ����	�Øϛ0��8g��cѼ��߉�^'�~o+��ߏ����q*�g��p=�T'��m7c����z��>���j��C��Z�=a#���p~��r����쀘�8=X�;�w��<�?��w?޸�Og�|j9��V�W�2���{����n��o����6��<����g��3��D�:g����{0ȍnNrJ����i=�3�4�����/E�4T��DFX��W�K�i��,=����?Y�Q���7�L� "��KwP2r�j�!]8�K}���J�<��?�RXT�[������*�J�t���'~J���g�,<<y�w�d�hu�QU�0��Lo	�}�c��ް?�[�}7������y�hS@m�ۏD6<���@O[v�ymk�	oS�{-f,"���09	H�m��y+�$8�<g�M�=�w�ԃ�Y`��,���b��#F& �������7]A �r�)��C�w�Y���\��Y&d	i[H,�<�%?���-�V��G�D�&KW`d�J��#�AG���S�95c)��\AN�� S_ƲnQ�=}@mYᝧ���s
��l���@��?F:��NXl
j�4��(}��8�,�{\_,?�:B��^�!��9Y�%n�&���l�.��J"B�7z\C0^���F�_�kŕ��FE�ĝ��RJ��\���a�Q
����D>�-ҩ�L�i�_hˀ�/��(�A:)�)2�d{�&�(��F�PJ�7�$� �V����i@���0gTҢ>�Tj���o���qC��O�ŬDICJ��2`Ѡ��@��w��>G��>���N4)�4�0�ɩ��ms?ڍ��m��ٙg��c|b����ԙ���	��0�݈�^z&nܺN�t*�c|г��^:�i8,p��O�w�'ơ}:8;f?�p�����ٵ�D���xl&�7B�RO�݊��I`G�y����i7�ש�~��)����,�]�. 8��zƩ��k��O�^�_%�Z̈s���k*�\E������|���E�cY����;|)�G��t2_g�.��0�Fa��	�2�<�a���`Լ/��B���2�������w�9�N�)��-���\
�Z����8|�:�����ooǘ�)>s�>N�Hr�?:�[z����p�7�q;����+����A�1	�ۃhL1pΎ���	7�`O8EF!n2p/�`��|�49�	k5d ��"��6/C99=��i(#�.lU�lZ�'���8f����E�&M�3kM�Qh�ǝl�x����?��v�_:���/eCdN���]<���&��7Ky��Bw%��2��:�]n'%,�T�����hV��~�&�X<�Y-A�?5.w!�B���	eJ�e���0�%<�,˖�G���%�$�"A*`����7��E��VI^�j#l���X���n_
�V{��:ՓB<S����yg}���`q�&�G� P��%ZAb�U�7**��l�ax��_�l��P�S�Y8���Y7��)�CH� ����p�'�܋�0�e��2�0�~4���Դ/�ɬIX��e���&��Єa�0��-u���y��x�r��!����C�"��TRcm���{1��c�HC����T��=��ggSi|n�z�����/Oh�\�W$
��ﶥ�d�r�A�P
G�$?�lc֣"�n{.��^�>���t�*�hu��` N ��B��Q�iW�"�V���|7Z7�D\����w����-0}:$��O�2�mi	���#��C��&�x��tl'��[����&7a��bmB�.�c���t���V�t�H��Т(�������^!�/�� YVϏc�I'��$0��qF�uU��m-x��\�5�t�/y�Es�K�RIS��ǰ#QTn�ԙ3h�A�����f��^;�,��!|ދ�?B����D�t�(MߐF�k)�`B��ƪ�:zZ`-��<��t.�/��P)�!��cx
���bo�x�_N�QV2\�£�a�6�b*G�)�&��/����<+\�6�h�f���Ϡ�2K�h�Ӛ��lsYn��tj�f����K����ٴ���;Hyfp{.��D���]
���o�@m��ya�WA�Xo2T5]�#���N$���P���H&����#a���A崪����}�>��z&$<��r��D*�m{��������:DY턥�>½嚪�+\� ��E#)|��9-���ڏ�n~a7֢<%]B�l��I9l.l��d\eP:�Hd�<����ξ�p�0,�٫���L�w���V`d����%����8�l\�a
���ifM�F�d>p�w����T(+�^�s7
ܾ��z4��2�hhya�� �$Io�N�a��j*��2��:]K�Rc���DwxP��8��vl�7��L�U�#�F�k0Ͽ�E���قop|�g�g���V��}���J�cbrKn����ܺ��˔��o�;&RkBѼ�-K�s�[�ŕL؝�	g҂4!p�Z�D���9UM��xt���ǿ��1�ڢ�����,���a(�x@	�:��������@��@,kQ<��@d��V���9��k��2�)�s�7\��2n��B��Rq�X��f�W	��I>~�3a��O~��3�R�iP�!?�/
+�� ����'�yTGR~���hlj� :��� �{5�����`)c���h���q|�w�w��4�q���4��q�� R[Rk��,�̽d��MR}v	p����w|d�X���~���P���2�'��q����-���^�y"�ւ$	N�ɟ;����|�h�t׻����+���|�V�T�^:V���rv��9F;���2ql�R�%��ڱ�?H/l��U��ց��H\�7��݆�Fx�<8	��TE�;Z��~f;iOj2��%%A]����9��k�ѷ���:w�%��m5�K;i�����&.�Rh��t~��)��۴�>%o~�����]L)\���I(>�o��9����|B��X���\�����uT�w�O!q/-�h��L�y��dx�q2.�J�@��va���|u���їݩ��h���Ґ6��|��e�X(�$�*In�n㻀:ͳ~��E
Y���ĭ�s#�G�s��
�k���9ʾJ�M®�{���:p���P;h�@٤��K�x�;��4��B�e`Ѕ/�}�b��.qf+!<��o�x��t��ƢtIW�/��娴V�{�_�ŉk��2	dNk�վ�. �]-^ũ�����<���K�MQ�gI�����/���8�X�t��J[Z�7֊v�E����Ok�|�gXS���G:<��O]�����e��3ۗA�lj�(�R�O���=?�}��]�kqI�F��ny�f1�F�ߍ����-4'��z��:����q�9�� c<�8Ś@X���i5��;5҆0ڭv�Oq��p�&�9�H�&�@9܌��kq��k����Տ����b�Y�S:�Ղ� ��-XHKB�����D�D��R������!a�H���h�N�rs
��i�S�X�p�	�xP�,Mt�Z���0�H��$S���ຒ����FC�}?b\�O��D�Sc����q�t"�� ��	�;)8��d���w!\��/D�ڲ���4�I�GؓYRt2Pˤ�d�<g�XS��K�#��As�x? ��7
z����^W�,	L� �NF��l�Z���@g�Ϥ�E��W������,����2�",��d^���k�V��Yll���qyY
i1�''[�
ހ}��:F[;9E��nJ��/[*�%̴�6&Sp)���nSW4���Q����]z��jp�x12Yj��0�%Mp��^��\O%g?�Ϲ�TLJ���Ǿ���,��gF~�zo?\.��r��<~9�xI�#�(܄QNNY@n^h���1Mz ��Å'�1:��Ͼ�PR���Z���F���%Fe!3>�g�U�q��J\Y��-3�'a��7�#nc���("lë<+rr��<=��9��&d�����7���}����%����}!a��ޙ	q�������z�~M�#�p�)��ÿ�T�\�9ͦ%�c�O�[��8:�s�9��8׈kK˱x�7��;���	*?v���H
Jzn�+P���˱nct�#_�F���ؒ^�7\�'MnI��4>��<>��M���,ƈS�(�����Ҽ@Ӑ1��Fsҏɹ�m/��7���c�d!��`�_tC��b�W;8�ڙ� �4���s�U�m*�]���}�����y{z�w��;�:z?f�B���b8�g���i7L�F�4�H�(`��_�0Oxd��.�?:ٍ�����E�5�!:_wD)e�Y�ڏZT�iU^�n;�/��S+xy\���S7O�c��~� t��'s�؄?�-ezkٌR�t��J�.��U�&��!��®�ǋ��ɲ(�>Y�a�_>нҮ�;�}��0m�B�����<���028�(�Ortđ]kP������ě �n��bh>�^� ,�����(�QA��H���)�͟��)�q||�
Yu֋��XZ�ʝ[�=�K��ns4>w%�}ĵ�
u�<�-�*L⹂�1R�SR�)j��{pP�'Sx�NX��W���)�]�J��Jr��|��~j3f��ny�&�(�T��c���s�'?������\4<Xtn��Y|�8�)qi�,c�,�hm%bq9�:X,*p�;Ф�z��U�_Y�Lʚ��>e�|�ZY#Ϲ�Nyď!�Tt��\�h�A�)|j�6�#�����{m-a=!�O�����$�������	z�W�BV��e�n�S
PŇJ����~T ��i(%�4���{�Y�����l���#J��YiM�ONu�����Ѧ���X�^����>������L�DS�3��H�6�hۧKe�J7@�ɰ�1�4g!J�tWn3�"�y�D�(��J�����i�[�
�%]�Dod�~7~�T��>�ǆ#t(0?%J^��q��<��,�Υr�po��}�"���T�~@ev^L P�S�4�Ր�4Z�>�\:���d'�a��6I�А"�[���k�-�뗠2H)���{q��v4�o��`n�*q5��'���#_Tk�*��D����φd��������I�n��G�3��(��119��U�Q0X8�]i���oI�% �2�i+�dN#v��h�=�>e�a
��ZD�Y����5�V�Y3&5kw11&N֣�{�Q\��6���((Z�}���4�Fh�\�eנ�uux��{����o�m���2��6�RhSF=���*\}����|I=��)N�L���j�+oȻ��mӰ��)��@aw-��2X���]q-�L'��$���jh:%ao�$�x�)3�κ�_՘}�S~(�*^��R{x��ũl��e�g�w*�t���-�
��,�VEM��ᚰ���G.���M��B�z�Hu��xw��ɺ(���!��ҕk1}�f��_�;ZS~-��1��>y�4�P\��z�0uI\�p�G�rc���i��`t;Х�Ʉ���Z��oc�&Z��K:�g��`׆��F�lJٍI@T#G!�O�3��<�R�G��7k������Bk9�=;�x�n�tLWy��V��2���=x=^���q�]^�Chx��,������=�/��\��'d�U]��g��p�g���fP��2z*�+g�$kO����R^f���V�>.c�P�.��*��岌��v;w�լ������*M-����<B��y��>C�a�2o�8�u��yIž�-cq����' ��g�y��1q��bl�V�nq@�|{�h�~��>�Fpq��Wc8���J���|\�iN�c|f�z&��܍�i��c�B��
:'-H��}�������@-�>W�����c;?=�R�Cx��� f��ty�����k�}P�
]����7�q�<ߋ��wc���{-Z���ۃ ��4q ���?���PX��X"s�6�?�1,���q�܎���8y��Es���������%ʝR�!׌�B��\�%>�$@�)t��OXI��b]��v�ύh�n�w��S�]�Ѵ�T�3~?�GY��3,�s���R�V�	u�#�m�����������Y�y��(Y?eA�*N=����^���	�
��kC�5鼗I�]�Y�o4���P��!�2Vj̫�=��_�d^�&�3�<[N2�,�t��	0�aZ~�C���P���U+빉��}G?��a���1<#��L� "��E2���:Cp���!�=��#��$����������g��C�.Ggf�h&�N���O�����t��3cp�<I�f�fNͧhk� �}v�g@���D$�ȓ�S+�t�ʙ)@��;Q��G�	�2TNN=�2-|�~���q�27T-L����c�#7l���"\�)����=�)a��'����~�=����bw�Wc{�Mx�.�OJ�8�O���(H��q\U&�H/^S0��+�@'wURQYyӔ�I�YXI����ql|�|̱�Ү^�+�t�n����>���O�T�J��%��4?�x?�G�|oE^v.wrQ�cBԦ���� �C�����ӆӘ�X</Do|	�ﴔZ�@�f(�d�	�M�S�'Q��(l�O~`��d�I��MEs�z��"v��h�B���������-�Ze����l;N�G�!��h�ȭ��D�_��������t,.-D���)e[����2�Ғ�^MU�Q�2��ܝ#M���Y�N�b~��_x<����S�����̯�9��<�WeZ�vA���������x���;�?{/N��E[= .Xg�SU`M�J
�X]u�M���}rM����瘖F
Xb%��I�������lt��т�Lc}�:�6ȟ���@��B��5��V�����|F?y��0��a����C���<����	����t�Swg������)G�)y)0S҃?I�0�Pγ{%�q��d�
���Ȳ��ȣ��Z���-��a2�"�l�!C��M��ԋu����|�%���sÅ���>�L�l����.UA�ӫ�0�^�4��9��`zǣ�8?U�G�����~%�/]�����~gfs�^��V�0���)|O�Z�Նֹvx�
9���B�Y����^ꗗ١y��U҆���@�6}5<(����&�[h�68-�ƌ�!��^�:W��r��/j%���n;�fs�&'�+8E���t���p��OaD��ɤ�����/���v��R0޻�i�],@��2�l]V@��_�D�g�[���H�Ġ��O\Y������O�&�m�v)_�$8ᧂ��w���bM�%��'	c
�j@xi~񋯾�΃���o܉��#
pͣT�P�b�0Qd�#��}Vظ#��n1Y�u��k2Bax�(�LaT�ﮗ4��jδ Ӑ�A�F��`y�0�;(L��	m�A��C��`Ne'�v6j�uu���+1�^��f��>�YS܄�n�-����I�B���ALg���g!+�����k�h���Bt�n��R��zJ�[>oǀOk�'�̺m@���Bg���l`<g�`� kwn1fW��M.��)������,�<B)���m*�2�gmH2B\���	������1�:7OVn�9빚!���ĉ}�ZaE���mK�3�7�x�1�ę/�(���6�e�ӌ�.JM����ݒ��)̬7:M!���ft~V�}�y���IN�Y>W��}"-�'H	OjO������~�6h%N�T<�	+m��m�����e�-���Ӝ�����)N�(���j@*��F���9;p�t�) a�E)a�����C�&��|�w�A�rw�̙��²����=��x�dޥ�*e���w��0����nJ�]��$��i�8<��Vcim9�N����D�d/F�J��i%c|y!FX}��4��$�ȏp͑/�Cw��\S:? Ͱ��!c�/ �EO+̶�?7�X���\�j�O�"j�u|]�lJ���u����f{����Opg�_�XK�!��J�J�ߔ^Hk��=��eL6���������x�@;7ۍ�˗b�굸r��X^y&N���Y~�1�q�R���&��g�Yt��o��.ȂԄ�_:$�fǃI�a�D*�c,�:J�P����L�_\{�z���.���� �"t
�K������{�?���q��D���=�>%�_��XW2`�u6�ѥ�,��y���c#Q�!`��ਝ�\�v�cM�0s���}�)���8�J~�����*�.e�`f#�Z�#0i�\q.<5�u�ǩ�/�.몜Y��Mx�,��7���E�B�=6э��y�"�j:�z-,Y6ɒ��O�˟�mS��r3���Jm�p��������hͬE�9'�0(�i��'D�E�ȗ0z�s�$��p�HUa�"�y��W&ҝ�6�a��Gbj�:����ˉ���C_=�[i��w�&��K��~�MҒ0�oן�:O��㳳899�����V��	��d?FG�[��\7"�׹��cG{�8ޏ����ʜ+���	�n2`�N�K�9�����<�hI�
sA )�V�6)*\�R�ʾ�Vgۥ�S�ݢ�(b2�,�X��=��r�2f8��+���|����:_�W@)|]�v86��r��Qҕ>QY�w7	_�Bʗ���u�.�'%Y���ZnD��==Ӊ�ř��x�,v<maHЇ�#��r�@�E.N��4���6Ǒ��Co%m����~4��rjn0I�)h���s���f#��YR�@3�\n;yg�ߎ��혞����y���Obr�oM�����Vv6����BX�a��;*�;ڜH(.�k��ձ�_)�&#���׌�i����E�e�n<>A���M�3�6��"�Y�(�P�J��J����^������c2M)�.˻�I_ڐT���E�E������`8\R���V@��C<�c$x�����{���?_��o2�Ѧ�M�6�������hUħ��r���֏ȷz��ܚk�լMa a:�LdY�\t����F��Zq&U/���I�	_nɛex�u�-xMoL���xK���<R��k
��[�h\��'�G�6(��ɩ6-�%��j�|i�tP3 Gj�N�h��ڒB^�$LP`�/A-���\8���;@�O~/�M:��P�vp6�hxg�)opJc�-�ZSp	�ET
@pV� ͵��H��F(�~�X�6��¼�e�LO�vx��#���i�����?����̴����$��)�ї�Qv��VL�8h�q| #���B<�9-������4��H�mE���-��)��鈩<Vb���R(t��� w4�ջ5v�N��p�yo��QC�K�Z��3�{��~�&Z��*S�8�sЪI�2�G�L@�S�.L��@���8�ie�R����C��,ˌ,�ͯ���p{�_B���5!��o%�=��0%��<�&�I���վ�c���-��d���p����ӓ�X�k�)��ً���mG�ӟ�X2��kf�_����$���z�P� ��}cg3ƾz�4���\��ш�Օ��eg��N��0߯��~�A���������;�����?SW?'��8����OF�Dq��_fg��h3m+��	~i�dhh�w}/�J(��)�H��p�-�'�ɱ	�R���:�7�\+�"g_9��G�z��az��: }ε�\fVe)��^�U~���O������eXU�<�w2GǇ1�ًa���j�M�ܥ,ǒ�Vbq�f|֎�O��/���6��q��P��iZ\e&a��O$�n���%��`+�%�����`�[�mNN����NO�)N>x��̗^��u��M=���/3��y%\�W8-\Ilj�i�_�����3�/�>dy�(|��p�QV���|�� $-edz�&iNW�_�0�Ї,?�-�����E}E�/y/�4�4�	���8f�:�o2K���ɦ��ԌK�JN�,0���5	��5��$�;�51?,Xz��k!�GhK�
5k��i���
 H|�G����h ��BӇM��vs�����8�xC|la���-c�x� �<)��ޖ)��CX�[\�By~�	;��Gc>���mFck=�7w�q�p�,-lO�M���f����6�H�j��a�2ڴ�mx˩\M�vUb���`6h��t�[��~+�h�-�0�ePJJ��V��9�M99����}d��*���2b�DB��+�F�Z��$�z��0�|!��S����oVb���T�@���1�u}��T�V�B��/�(<����8|��G��;�'
ĩTB_	'�3\���C1�}�9R���P�"Ң�a�C�C�&�ѣo)����9O�b�6Sɡ,_���"���a��D�qKkϠ{\�6J��|7�8t�z(�?h�c21�@N�f[K���1�.�D8y��q��Sy�4��F�"Oh�Q���s�o,4��j�.���<��򍺨��{+�ǐxn�$����7����72�r��1ݓzs��E04��q�����1��Mh$��Sg���e|F��T�O��^���N��o?��C�ZS0R���p��8:�&���+�y��0���&���b�O"ə's���p�>M8�N�5-�Mo:1�s !lFY���"�����&Á!��S��4U��,��6���KS�s,Uޒ��0�/�cfB��8��������=��M�A��t�&����Ԣ�TN���b�[~-˭�
iaɾ�O�/wJ�D�nK��JOp���zN�p넳j�I��ܦ!���[���37��Qj3�Q{h�*�Y���iɹU�O�<˳bp�U�i�}�'q�G#��V&��ܝ����}Ç"ޏ�}��.���" ��Q�)�V4�`����V,�N�D����I?�҉.�u|m2�:q�^f .�ë�ۣ������0F��@��BwJ��8��ќ�6�N���噾�/���st�P��X��^�P�*�sי���з�����d�]��3 �����l�x�>�S�'��.�]�/λd�����t)���N|�K1<=F�	ڨ�;X�%��:0i�mъ+�,}*|V`h�:O�	�aBN_������TO�����=ދ��>�zB�
}�NL���p~�`�	�]����&Y�wt|�G��x/��{�P���x�Wʝ�b|�C��ϢGib�0<2fbr>�^"��蝷���<OWҖ����c�{�\�R�{���9Ĥg���7.�e:~�������ű��E�w�Iu�~"H�}g�	C�	�d������.+-tZ^���4�3��*�}��-'3q�gpl9֒�������%���OW���[�mS�s��oa��D�5Pd�
�o!|��}:������"�)>Z>�p��!V��U�6���Mu��$�M�H!&��}��K���CS�_�RE1�!|.\����:���ag�R��E/�[_e�����'��4�Nǵ�Y�p����RQi���f�$ۖ
.��f��x����i�%�(�th�ZjN0XHxR��:$�,�$t6>�=˲x��SmnM�zq">j)��K�N��D:�|��i�;�q����iNcƜ���d��mqO��$qN��"K���hN�x ��=B�و������C�p�6%,D̯�cu�W(W��Ύ���F\�jĥ��X�8���^,M�YC�Xܜm��K�x~u:^�2��X��k�ѻ6���(���C�a3�z�1�D(1�|A�C��сS��V��'�w���>�Sʟ��;VH�x��m[|�:�YW�tV��ii��<���#��&_���a%"���i�,W�N<���-��>�M��/p�m�)�ssi*�-N���Q<�9�C��E}�o��mz�t#����:J��dT�;/S���L�#hˍ9\~z�X�m�"��$F��9u�;+�s'����3��Å9"&`;��)��u�`�,�!V�6x��}������A�K[��>[�1>OZwP��Ɏw��f�VK�4>��5��d �N|'��>ҭ���g�#�(�L�Cynؠ��������F"�W��5?����ٚ�X�|p����8�����x_+��[i��\�P�BK%G8T�Z�MO����~�2�J8���9}�X�i�I�9����Ы_۝D��k�*�YE�f���Ռz�p���G��[w�/�'�_[g�S<���EN��)�-�10>�bd�4af	�]�'��{�SC���8��]�t��
{��y����zIU�qYC�L�o@�S�9���_�:M�La2���+B3M!A�%�	'M��5�t���:���$�4*�R6��,�{�>���ܦ�N��L������:2����-�ȧ˦LۓB��$s
��9�͵����v�h;Q|�N 7�K�NǙ���2er��怲\�&�� ]a�֥��4�Qm,���H߃j�+x6c�ǵw@AZ������XX���s���.�T- @忧�|�U�F��+�l�4h5NDk��q,�I�ec�Xµd�c�׋���x��N���z����K�'vl� �]����ז0,���ŕ���h�%�9�@`Z�<�)��x�9U��4ބ���Ǩ����;/�n���WlN�ƛ[��/�)�JG[~aV�ɥo�c� ����A@H�-���Z�S�-~�ε>S�p� ��š�i�����œ��-,`����'=��H4y��s�����ٍ�=g��t�Tn��e���T�⭇�X��ฏ����a-?�C1z�&�FJ��c^4����c������g�1�F(��1��	.�93/-���k�h�E�5�A�XE���W@L���ˣ3��&­hөxiu��q#թS{Ԓ�����Ŀ��C�C�����N���v�A����'��If�L��QI
k#�$
�Cqu�ˌ���*��M��+H &M}^`�@p<_�ɪ*>%��\�	g:в''1~t�K29}~���ԥ3Ίȇ�]ɐ�3�t�����_��#6���.��t��X���z�T���&4�m1�Ā��|R�Mw� ��ݵ"���㲳2	���p�I9�\�MxIo��A�M+�K�P�Rqc�V�&��R�������~wÜ9����RJ��$u8�Q'�	5]i�Ҿ��g�'�!O9�� ��	򦍖c�[�A�Y� $�����\�)�;J��,�G[)1'C���s~"�r�2pY�ږ7���#Ť����Z��!�R��4�s�N��5L]�M��r�BV��~5\�b�9��
��pi�j�]{�����O<~Z��mE{�+˓���2;:�.�C� ��{�'C��Eq{�P��B�mu:љ��Nw::����R0�Պ�n��,6���-��o>��7ߋ�ΛY�0������b�����D�.*M����8��M��a��D��	NՌ�xI�O�`�v�|�����h�<c��G����$����Z�q(0`_���Oi�R�[��1�IW��x� Y�}��O���<2�9�3��q*zI��+t	��Eb�S䴚t�H�����X� Oމ���fln�!L/Gs�j�ZSqr.�S9�j�>��w������f%��c��1���⣟�(J�Y�����h�0Q�ks1ә�������3�o�ǟ�w��h��_AO�#���5J|�>ZF��D<s&4���l� �t8��=幇Z���D�C_���k(5(��a��א��shKuTܤ2)��K��ݞ��P����*�cD:Fh��3ױ<�sZ��<�O��h���mv���Z����*g~��֬�j7Z�a*�&y�y�<S�<�8c��j��"]Rg���Ty��Ǔ	}����V�>h�1W���'��������ѲF��߉���~36g+������~ў;v�7cr�a�4�(X$�Kll�'�+�1`ЈE���--cF�'$Ȝ�/�s����]�dDV�x�c��00��'gh)2N4�4I�=���SrJB�2��Jd{�ΰZb�v��ՃZ�-�:��	n�Q��$�8hOqXO�a�,��Le�ɼ������3�ZT���&�t6�["Ѡ��MR�6�$[
��,;롟Z��3i�J�D/�I�Sם�T�
=���+��gA��}I�+Oώbt����1���%MF&97󳭸�ԉ�	��>	�/�a�����
g�h������ �VNgj:�g`ZS �/�:%�[��K��Yj��4��N���n�v{#���o������i�
�!�מ��U��iyǆ�B�qï��I��YOU�$�#@����c���N���=�y�qL?��Ѽ���Y��0���f�c���]>��E_�RqJ��fr�[rE��-�Nۗ�a+R7��LN�(��1��&N��uf��0՞@�c�.B^?!�0=���qp���~�`i�Ek�V4����\��#a�����K���u��x�������Oĕ�Q̌��dw'޻�ocIm�Tw"��|&��/���B��'?�	ʃ����)����/ǿ���c�~�?�.G� �ӥ4�y�� ������
:��
�+yə39�T6�7&����=h?��*�%��K�K��X�Ed���T:�)�<��tH�&�B�5�3���(�%���W�y���w�N�dv&�����G:-Ep�қ$?C���PeX6�/S0�l+����-�!h�7o��`�����8�!�i���z����L��T�,g����
s��|m�H��Pb�_��^}��A�̷���wAlp�d�j��q��S�`ſ1y��ւ�#�fN�q��j�-�?0�ìv������̸~��+8��,ý��y]L���6�D�F���@8�Y/��g�+L	�0#S�볙K��ו6��'������RV��/�|�,V@UV���D�7<�e�JJ���p�d�Py�NfQz��kHںŢ�WW�ʲs0I!�1<Ӌ�R���e��$�lWV�U�%��L'���(~J��AK���n�&��
`4cXT�u�;�����5?��8����-Fn��Ҧ���q�6v�Ok2��NL"d�S��N#x�z�gfc!455���:\'�XE]�vq~1֖W����x�֕x奵8�z%6{�q���<�n4vbt����^߿?N4(�QАE955F��w�`2!(��&=��[G��m�����c��+1�t3F������C\7q�>��(Y��}�k�\�:`����7��r�����? �}|alSL~]&��~s���=�F��w�)�����R3���;�����x�~frK�pi)�V��#�8>-�_2ӓ^Ll�KO�����/�����X|+e{�nܻ�.V���;�A���C��+���l;^y��1�eX�4�$�*�{�Z��ݯ�7��u�V�}1�n����$H��u�������9�QB3]us�	<��(1G_���j��LK�וa�௱\ƌ|G��]�e����)�$��S��x(�	,A�gkx2�:7�do�{�D�%�����*p'�e<O���gx�G���>B�P��Ә�I\Yå�)�R>��5ᾪ��5�ทz��慩�1J�^��<Dir9ƌIQ
�g$��k�Z�~��W_}o�0��������'#���Е�#�TЖ);�f�X�E���Oi�dg%�e���+�O@�����E�d%:���<��K�?�E�eޓ���wz!kW%r�0jA�����
>�r+3�(c�T�z�T�w�����[	�t�H-S�ۺ�p�c���HAT���f���2�P�Ѵ� �
�������ʴ��H��?ɭ3�ɕ:�7��lx�xc�s���˨)>�m�����T�ӣ�'���Ny�@��],�G��F�G���q1��{ӳ%ǎcn���1)�"q�G�HHV�}�֎S�-���ȗ�(�13��S	�����M��j���<7� "~�4=��cSn\��߸�ܺ'ݕ��a��Cpp} �FY��b!�J�Ǻb�k����,��K��0�@F�sS�Sn��X�������.Z���0́���}Yp..�{骐Y��/��œ�&3kюɥ���pt��lM��"�O��<@ؼ�ɉx��L�Z��9ؾQFBY�(x��4C�N��Fi<�r삓g�6֮_�����q)|��r�P'H�[��G���~|9O�_�|=^����S?�����>J�&bzv.V._��k�c��-b�6�Z������o�w_\�>���v�ma%-�t|��b�ƣ���%��\GuV����@JZ=e�&��.�Sm�n����K���]fs��7}�+�����~������$s����X�q�ϸ��z�/��;(mZ��C�/Rcy��a�1�ܣ}L~�Ax
���� q(	}���~���39yd�<�@:��O�A���g��o�Ix���S���$X�h�A1����o?܍����q�	�0�u���d�43�
n-,�-W|13�;��ܞ��̊z��3�*�b��L4Ԥq@x�,��c��?�������	�b�0��b �{0�3�O�<����G��+5�|��i��[a�!����r'�/\
�tU^\�A�϶���3&��+!�6�E�wy%��{)�t<f x��.*�}�D��ӕz��P�Z��>G�u.�ƄO��>'�#l���%�b�Q���T��hnd0��ÿ&1H�x6�! �s�4�V�<׈[X?����%�/��IB��?�����O�8�8
�.B��ʙ-V�֏qm�{�n�2�N�թ�.iLn'�>'aX]��<����j��z��R4�V���i�l�\�0 �JO~�2p݊=�� E�f䁺е�-����K1�n��e�V��t4�֢9w=NF�8��?��S���:�z���O�)�����ā����f#�F �[�(_��������G0������//�g>t=�C �3�wN:I�ٷ9�y�@۟��sњ��c�՝�K�o���l��>�����B~��[0I?-^�:����$~�c7sJ����}r��31���1ә*���]-��\3��wߍ�?�c��&�h�l
D�e[T�NrW��	V���"�}��ꌂH�U($�f��/��&2�� �_���|�����ȓK E+%� ��jao����K�m�˃]�|q�s�}�vɳ3ݧ�=�b��A�x�8����,C~���S�FI?�{!N�#�/�墶��l�c2鐫�0F�S��`Qf��(M+�����.�i�D�/ዯ�E�~�w���# �d�{��%QhS�up���`�&���!�y��&����9M���z�v%���P��ct�A}�+��������ͣ�DcZ?��C����h���p�h'����V�ʈ�G�>��:>�$���AP�ͻ��X�ė?��'�0f�_�uɰ�dc���#&���%��+�d��*���Yj�[�L^�+���ܦ��kkK��ė|UhI��V�Wާ�ZR�2?D�0�Z�ĒV��t�����ǧ�1���<��7���3���ч0�5�O̢q����x\�F&�i��\0��PW(ؽH%���! ,�9<�n�]X�תq�L�gzF�3S\,�73���ʵ�J�'ׂ&Z0��\��9�=��7�g�c���7֖cF��;�X@C���N�i�#��ږc�1����;H���Ң?8��qK�1��4��bL0>��:Т�1�^=�+�->�A5�
�+�/��Y��)�IUx�s3Iz����Ƣ;ޏ���?~���-�JX''�,��E�����q�&^�E]�[��S��Ķ[(��q�o���~��?C�:���8G+G��H�|�C,������>z5��i�eѥ�Ζ��6JCn����4�i�g���~)~���� ؿKD�!x@Ev���y<�;��c�9Gx�բ���n�u�F,gV�[	ω�d�^T�[���8ԛ����;hd�T�8�o^���,@ `�nE����]��>q'���D�i44��/�W�ؠ��1rNϴ�${�=���\	8��TU�r��	+��	��&���3��Oe޶:J�X<��t?�h9u��KZ}���r�ZL��^%|����|`����C��vJ8�窼0��\�+�a0�Z����=G?L�>����6��2��5��e��wv�qp�t9jɾ�QJ�Oqa%6�� �����<�:����}D�m���)e� ����4�l<��,��t�^��D���XI��<X�s��򩘝�3J�"q����fRJ���/���B���/�k�!�ʎ�TC+�a:��`ڬ��'���t	�7�-g&S矮�f^˭j,ɹ�^(I�M\�x �9����X<�1��_��J3n,O�U�(��~6؍��f�uS>�M_PxsL�&��^[=����)O^���So�
r*��.��"xf��"�d�%7$r��S�t�)�ܚh���t\]Y��gc���Cٻ��	���HA� �����A����4��Q��,�gZ��mnn&��<+o�=Ð�r۶���e���8�/�yo�ɲ33.����[�j�~2Ó*Z�:�F�����Ka^Ҵ���0���q��`��7���~>�Щ��b�����i�'y[ȗ3�΄��2��a4�6a����A|�Ǟ���ZZ>�yw2:A�S%���xq����W�Ui����_�_�{�G�
x��1��
�G/�}�`��b�>�;}}o��
�U�kP}��d�S��+�3�����(�R��SV���s������������L��bm�J��"�E�[<Û}�{�^P��Z�{$�p�{��c�wk�Qy��!� �x�˺�!�!/�������\�g�����#@]��/�_��6g�ɔ�&uI^�(��ο��W߼��[�S	�}D����	���-�)�:�C^#����ĭ&�å��l��|�q����C��� %�.!��up��E��%̶���A�!��j ��#G���D,0&�{�H�hV�w�=!*#J���՝-�j�2m�����D%�T���,�rK��C�땐W��SJ͇ߛ��os�/o����Ģ�-Wpy2��/�U-����T�Z���Z`��s^��m�`<~���b�Q7��뭸97���X�G�EoN"@���� ��Bf��	`�cM����"�Z�)�ھã� i#X�0N�9��ѭ����1�"-��'Zs 	{A��W	�v�6�ø�"&��X�����+��>��"�
�'`tX`�Rc"�	=�4JS��c�|�@������S����qt�[�Ք����.?�b��ex>V�Ȇ���\�0T}*�u�J8�s��c|�n<��G��"^��\���U���x�p=Ucc��&!����1�A��8<�K�Cs��b��:Ȗ�)p|�10n�D�h1>�#��}Ꙙ�
��70����U�_��Y��/W�t������k_�R���~���<�>��h�]�-�$�'$���O���X �d���JH���>���O�=i��
��
�����JJ]�3�K�3��.gg:ی��(��O��P��8��_�o-���tt.�c�R+f�����Q,�cy�,V�.^j��=2w(3�[A6v�ng����=w:���^?��g�����IS��/}���������<�Ϟ�ivת����o����m�G������{����u7z��J�	��8B ��0�܂���/LI����Nw��3
d6vb���� ����׃JՄ.���1�,��F�X�<���{�h�y߇�281��@����$۳q�"��>:�>�T: ��)E�S��E�℥z����ǫx4�����x~�%h��@_~}���+��`ϒ��M!�V'��)W��u��>g�����v4�ʻ�/�K��*.c�K8.�D��y�ϺܴP'#]n_�>{�̏�m���f��j�rV'���n\�m#|&b~�����X$��o���B
�jƱX&H�	���~�$w�yE��=^��\ĥ�)�]p
 �W���+#�Sr��v3��j�Q� ��p}k�<�@��X*��q�c�m�����ԉ���}9���S�sz�i+��Kw2^���XE;�?<����8@���_�M�N)tQ\�t�+���G_(�i��޾���
�i�3b �'�q�ԏ�u��c�ڵh�ۍ���>JH�K���X/0Y'��0�f���&k��d>
o�C�&���N�U3-�s�x!>����4�r�.Ɨ)�r��T���|'f;Xd�N�l;u�P���oǷ��[�����C�²�G��/.?%||5�?�.��Ɩ�-~cЋ���jM|�����"u��n�j�A�1Ѯ���8��D�]q��|p��Bȳ��a2�1����`,fQ�V^���?ЍO��j|���x��x<�Ҏ����،K������x��\<�����������֍��Q�� ��1j�V�$����]g@�J��sC��7�?i��!���(P�2�t�@�O5�"9?ђ�\�*���r���?$&��Z���_{/������
�	����RYl�Ҋk�!`:P���N=*���Tؤ�s�y�	5<�9˻��'�ݙh$�]i���ug+&�:���\ܼҍ�0�٩�o7.����}@#v�����ޏ�7c��N��i�֟�>I� �F�<n�sΘ�;��~jw�^(����QQ� :O�&��IJr �T�)�y�9~ĩFt��8wc9ϯ��k8ً��2�Հr:�:�W]*��C!bG@	/e$q{�_�/S��Jǒ Rr����!ьƜ�"���պ���Y��y2�va��mi�kꢴ�5�3�2v�B�����|1�PZ�ث�X�Չ�;�����0q�:�
�m�q4f���;���K�ϳ�/['�hծ!N��N��[9�ZQn>�I��7��\�A�aAu�W��M���W�U+m�I�|�Z�Ö�^�)���oo��/��k�W���"���/@��h�2��Kq>7�0�h�z=O<S�χηS~N����k�Ҷ/4jeh��R`�N*}.L�{O�4��=?y_����h�P$��:�k~��b�{d�#$|x}����x,/y�B'�aҏ�N������	K
+;e��@��в�(Wi$��?7�x�����~���D�e<��ч�3�������O����zS��hǊ���7��?��}�ftg]ӎ���[�����������/���c�1?>�l�ǯ��]���B�����#ڱ�%~��h������T�����L7����pڪ�s��~s�bNɊ;���-^������&�v��H���&CvH~�:��!�\�]Wr�4o�S�;R=����͙��2�3�Ю��i���{�O��0��&�7h�#�-�L��	�����D�9::�=��#�bq=�<�虊��Iy{s	FPW���sz�q�ɱ^�U�=4��1��=���
V�${��c�R��E �eg2~i[}����4�p�_x�����o�Ư�LR��Ә>�q,��� ��#��l��m��� �<��v�c��>VGc@�6LJD#��D��tw!V�㓟�~y>nݼמ}6���#Ձyr�Q��.3R��t���^lmmb����Q<�܊�nߍw߹��~l>܄At!�%rLC�Ӓ�4|�j����ԑ�f��|
��Γ�'~�+�s�`B�I��>�I)a`��J2�d܅(M�sN�0س3Ԯ���vge��N�aP6ΰ�T7�PS)ﱔdB��ڋ��n�ܗ3��?��d�V���s���/��KHl�^L9��؀A6:p�Z��ja��ڱ��ps����W�V�z>nD<�ˏlQ���\���^����}�ف6�D"���x ��5��I����%�kD^kaKiY��.?"<�+�+d� yҌ�SJd���G��_��W�?�+�E���/Co�h����1�V���y.m��d`�IE�9�G���Z��Q&�P�~4�� <��;R�`ִQÝ�L��SB"���L(Z�zSѐ�����l��8s�_E������L��/8 d�v���9�y���V߇�r����&�[���^�޼���u���ۀW�����տ�'�}�f,O+|�Qe]#�vl@G�{��q��L�ί���<%ۯ�~��;�?���7����� �l��Kp�Wb���clK�[^t�?�4��=��U��S
�٘^�����8$�B���*"��I��8I���>�V�3�����!>�S�e��[6X=>�ƁJ�*��
ߩZ�َ[/��g����JL����1��Ǫ>��b�{��!-cD@�N#G"\zǋ
�<��R��_�7���!�?>�w�o�;w�Ǎ�6��3x%yG�I��� T��{aUШ.���R��������!��AG�<�B�x�����S'���/~���{�^��w��Z{�NSA@�����|���-�4�↯�!`�G��V4O��0�6�aB״�ڱ�Ѝ�?�\�����������d��&>��q��J�y�E�� 끐�ܽ�Q����3����y��/={#^y������W��=,���=:a±�4���\s�ͩ �%-W�7A�{�ɫ��1�eHhe�� ���9�o��Hn<Xr���|R�q�ᄧr�yx�t`�+W,�5<���Y�7I�U�[��<I ���ĺ�?�.�� �W��*2�'�$X��s3A�8ƶ7�pQ>���i�h썙X�ų����-��RL�ScS�X�n�FkUP(0�S�p�5�;ֈ���Rs-�L������=���1�� ^�S��~�))i:�J�3��Dj�Z��� ��C�l�V���D�'�ww�����.7.��`���L�!Q	��O�Z~i�)�|�/�&���$A����V��5�s����oE���Є���Q��<A�gl���C=�����u��En�}�N�]Z}j���p�-ª|DJ��|4�a,_�H�λ�yH��]p����Ǐ���qM{��	nh�hh7���?;9����8�����VYc2��{���k�,�<�����z�~� ?9b3�N�e���R&Mh��_xn5�����I�d��������<���|�p�3״0�]�+��-<���_5vw����� F�0����$�O��J|��7�^��\[�)�n��0���Q�Ctt��ǒ��.
��B-��"�d�}����Ԁ��
@�����l\E	��Ǻ9����ޱ,��� q*j�9#�ܑ+�?��D	Zr����d��,��n;�r(�STT�K��?ޏ����8��IH%�y�I"U�h�������:@yΏS���Q4�iR�=�˯8E����\�����_��?���c���?�<{�n�>�j����z� �߽�`ۘ�Ǉ ��0�@���^�B��X9�6�����X����cum5V�7�^�+W/�)|x�ܯ���8ã���O�.ߚ�A)�:X3Hy���&
 �J�^,�C��<���Ħ3I}��0�Nez/x��p~J�.C*g~}����䟝��Ilҋ.�N��*��P���A�_��$*�>�f�L���SaֆRaj@*1�j�(
#��X�ߴ�oD��L\����X*Ͼp3n\���AFA�F�J!���In��}�3�f��5T
���3i�+�`�n�������yn�Y�/�Rn���KD⹿<�3��Ƨ�!�������A8	L�n瑩w@�nG����)�tc�Q{�<rE<Y��9CU��A�pM� �m�#�:����])���ʬܗ�L)Ô=_d B�5-/���〃a/�#ߔ��#@�L������y`��؇���C��&�7�j�'��M��wQ2���r0;;��f���r�0����L�LM��%�w���x?����w d*�䝋��c���3��{w�;��n�#�'��{�г�h,hQ���8v��6?d�p7�g��$n,n��>�{���+m�|���k�i�/�(#�ۗ���g��x\������~��!B�1{���R�ا��Ǟ[���9N�n�8��N���v���$��U�����I����N3N��fc�����	
��G��v'&c�ƏC��,�cg�8���^�'��>�0���������L�k4����Џ���α�F
>�����!D�L�ʋ"�y,��ߎ?�W�_y��I�z�\݃��Pf`�0T��8��(<��6�:M�| ����k�q�֕���§�O��O��kW��#�(�܉�w���JD�a�� �|<��O��h��mۭ6ȝ�X;1���)>���)�xp��i9:|���}_�����_�f<z�}��uz�q$@��5Z@���c��ٙ<ܯ3&3�h�Փ'�;����r�$R3�b0�֋�D��teg�!%u�E2�'a��"���AR'�+*��.��ROɩ�XJ��Gx*�C�	�� ��C��.;���F$V�������|F�U6Q<���H�v;!^n��k�����_����Z�rZ8���	�)���>��/�$	��(� �ΗE�ZK�@�>�@
$-����H�;O�i�)/[j�R;$��ub���/ָ�S��(f�	� �i�������|+�����w|��?�����G"n^��sʷh���A�ٗ�et��c��Fj�%�IW��,d��&в�$Ig2���ֶ'��H�����S�kɾ�EƊ��O[�(�eC��ժL*�$�1��W`��&c�C���d3�a1=���ø{i)���ǽ�8�8�m�XY���E����ti.>u�Z\Z����B
v�	<gkFy�E	LN)�ЄU�T���3��� ~��~)~�������7b��cn!6Y���I쿽��� �8��N?���[��:�l拶1.� ������#��u�+��1�?���A�ԁَ�!*q��x؎�=Η�n5\?��̇�ӟ�/�\F�f�����an>9GI��O끒-��X1;�Q^>�>j�O����?;��sSc��Y��{���10�b�nai>�Q�Az�B����[�ߎ�yg>����8?�<�xe����V�R��h�Sq��5���M;y�E皙k˙J�1�յM���\���n���b�wb�TnL� |�g��n=cđ����-�?DýH�� �c�97��Cz�F�s��G������3+K��?=9����}���s��	f�[�<��'�Y���i���h����[ggfgciy)��;�)���13;�Ҷ��{�o��n�������.o�_������Չƥ�hb�b�%�ج��"�Ɍ]�!`�ED���l����!�g�=,%>�<�2��� ����S)�ڳN���I��J_Ց�]�I���Ŵ[.!�',��g|2j�ЛZ�å��'�d����l#x|�ԗ�����y�o��<��s�~����[9��(�Ru��I��7l�mv�� L���w{�����/^��{9Y>^Woe��;}���]����sN�R������D^�})Q���������?�������?�Go?A���^���#,kW���"|D�t�U���bMZ��?i9Ô��'
����(�dɐn�q�!�t��C�\%�M�5_���l�}i��~�b��c�1ܧ/Q�TޕbZ����o}������k�h��{�Rq?�?�D��O}"�\Z�/�1ߙ�?���ͣ����:k�z ���Tk*ZmO�vHM��9���ȁՃnUt����y�rzڏ��8DH5�E3�؟v�<����[G�K����+��Wb�+�:�B�	J����y����iA�!8}C�����Ź_[���h	ȯ@�_n�r�G�r��p3��җ>-	���M����}�R���R��`}#���r�}|��/�t;��f+�orJ��T�X�F(ϩi�M���F��P�����~La�������X���G����{9.�f�c��j���w����>��(����<��s`���څ'�Kτ!���m����S�=�C5�Gnd���!뭼0K�~��������[�ݍӇt�[n�ô��Z �x�����q�A�y>T20:c�ڕ����c����L���a�?E�R�8�����o}7^{��x��;���8ΐ��H��<�a_�غ�����N2|�^��M�-n=#�	����'!<�v&aR�s+3��LO-�!Z���C�<'b-c�U⁊�|Ω�[@�L����<�qZ����4��U���c�L�M�̧D��<�<�����a1���e$x�"��:[�S�iʵ�K@�J@�8O=-�%6���/u@�$;��57��Q-�"a`0�Q��0¬����ћ7��4
Cnw�_���R54xZ���^�q�ZN����<��[�|��dj��X��NN�1��hu>���AYV�F�l�(`�3\�5�?ê�Uz���9˿ST�ߜ�j�7Mu``��͍�x�ZѮ��e�yT�t�K}i�Q�`ո7LI�S
W:1k2��ƃVh�p��P�>�28F��m�,��qc�օb�U%c���p���Q�[1�+Ƽ�-h��=<�tl��Cp���R[(p0{�{����_���T����6~⓯��_�������XŢ����/�.-���BN	-Lσ7�$Rffk���M@��5���n3���v7���\�V����h�af1Vbmy>V�Wce~����u:~�K�sq%uyq"vމ�~�+��sXw�6�����<-x�wtj����q�As�9�0"׿))�~s�{����h�s~-�wjm2~����7/a�cc�F#V����:S�0Վ9��4��!�-� �P�3�9[ছ.�2vƵt�p�����;��e��Tg:���f���|�2�
cm"P4H��q|�3����p4�xt��^*��eO��݌���s��ڹQ"�Tи%XOTE�ҭZl�/��/������[�{�[��T�Z>-v�J�Q����9R.�v��{�U��p$�D{!������8���O�󗗩X�3�`+��z|�_�o}�[�����a�� y1�s!�V�Ђ$�I���2� ���[�t7��i��Y� �@b�F)'���qkw?���v�;�Vf����q��6��l��!��j��@�3��@��[���A�QW�G��q�ˁ^�K&�����7U8�����xG�|���W�T�f�Օ
��M�.?�Mp�qu��t�j�2���Cq�.�3����>s�U��^!�6�蟤֜'x��k�S�h.0P:͸F~�#�g�߈����Ka�`A{˗[�[e��x�<��m�9���a`��qj�i�&�T�g�WD�^qV��Ҭ��+A�-�N�)�엪ٙV�R �֩Ǒ�M�<��!��J�f;z'g���>��ͽh� � Ǧ&+`�"����{�9��>�+��uP�t
�\�3�*=j�h��T�S�X=.K�w�(T& �u���f�NQ����p"�����e�����G��m��Ÿ�ƭ~1��[��������_�_�h|���,WŰH���~������Y��Wpyi��E������J�7�Ȱ(+q� ��v��Q�x���c�����W߉�4�x)�=%V?>��qx�0�zV���N�9��G�E�5���F;��~/�����}�%��vƱ������������ks���x��q�Сc1?ӊy�4O��-����sJΗ�'T���.�?,<��n���9�Ռ�0�M�P�L,����K
��1��^Z�J���`o�c
�`me-�K=�C��pD�{`U��5!�גt�r��:�k?
��,ޓ�	�l���a �����W�=ډ����8z|��"��z&
�B�i]�k>J��; �1!��w���ϼ����D�k�Q
�2�$0��Y���Ưǯ���o�o3�r�M�2�Μ.�a���X�TkE 4a0���8'%;e��C&��[l��_H̏�!�����H�3#C��S���V�� �; eg�q��t �@ ��)a�?��af��'� ��g0O�cD�D�S�����&�/�gD%��\���8)E�2�����j|^��8r+�y�#RF��׬�$.����q��c�m̺���2���.���2OF��:���t��������$���'Cf�2��K/���}��I^�B��~k�n�4a�����q���v�B�n8�`=� �j�YZ��+�
�l���^�/Vm�+����a�6�TYF��B�����YW��X�4�??�׶�c�,����|4��7�����
.n�#�R�۪R���%���]��@^߭�vU�rm�o���xP�54���������C�_�Q4Gj���i_z�u�
brSKh�ӴfK��c�ſ�/���W��?��Ǉ?8y>>��\�N�N	֑(M�%�� |��%s%����9��'�>)���6o��8S���fߩ�[D����x�^���ͫW����s�����ќ��w�z3X
�0�),�&4��H��U��w�h'�|i*�(*��]�<��Y?��c�=���X���?�#W�/.�d�4�?���7r�K�����$���Xth��m*6�a���9N|F~� @�Sj��'���nFNGO�d;&r���H+kh��x+�����ggbyy%VWW���+�l0�v�h0??G��8<ގ�^�e@{���2��`�i�>$��Ji�� w�';���ٗ�$��O����܏�������g
�m�������d�G��hD� Xkm��_����?�G^�Af!j�;;�㷿�����R<|�6�A�LN�t�ڳ���ٴP�f�X��EdT0��x<�؂DO)�����m!w@)�ܞ�N�1�I�bBMWK�O O�%���aI��O��r03����Qh�N����ܹ�}�W������z��螉G�^�eg����;,�.#��&C�շ�]2j�k&��E�gd�?U�Zj�*M�/vH�,9˷?)ZB������J��VZY}�e*�=G��`Z0�O>�\<���|q8�Y�/�vj�~�E��uȄ�@$�{N��7��2˩�*^�d�*��\���p�2s|u��m"���B��u=�+g�uiy_���.8OO��kw�p�O�F�(3
�u���������,��Q:�;/�o�)O�,귵�Kv	b�qw�;�Z����<�<��g�"`����9�Y�����xl ���t��s�S����H��?���'>��1��"���ԧ>?��Ob���Z��(�ڍ���S����.4�l���*�d��S�+��맴�.���U�ԥeʋ�+�}N�������wb��{��`/]���t#��-Ek���\\����~�'�?�#���+�톇��S�p�C�S(W3���{Z���|s��n4��5�����g���?�L|�#�� ����};�~��T��z\qGZZ8Y��n*^���Y��Uȥs�,ǂʸ�(f9V�/�#��F@�3U�I���˴���x�����ښ뛃,Q;N���>u�b�<�b��G�F�hxH.햎�v��V�*|r �X��!;���tң�&(�͟��O�zgc7��w����L�>���G�A���;T�9DI�d�Y�+��ޫ?���} �	B���x{#~�W�A��/�|<��n��I����� p.�c����	�|$�����8��s�ރl��~�cX��? �@�8lm`\�Tm�)7��e����s��t+�onގ�L�!�h7�/ܪ�.����Z@��)�9��ȹ:8��P��|6/�uP)�K�z��W��}�š��P �i��T)R��.��"�J��3��&#���B�W��tyr�Ǔ�]lT�k������o�X�?����ͫ15�@�Z��<�@n=.�\��
�S��spF>�����/���
�z�J��v����e=��=im���歞�/ӱ&{U0������������8�]�X06�F!��`�P]NQe%�	0�Ib.I#���tmb���LƼ��A����n�?�
�CX-���c���A���B]�M��9���ўSmЎ�>�B����?�������>�����}<~��X:/_��4��Ǐ��;�!�z�
k���('Ig �  :C��X]�h�<-�����D�S�!����o��'.+�pZXg��}����W��o<�5�׵����իq�����L���s�'~��O<>��t����ʯQ�2\�F�r5꺅���}���~�ܪ�t(x��6�nď�R�L�Ž;��{�o# �Kqii>OMGxi=h�IS���q"!H�0�^��A��.�L�̱��Q� T�X�_2�R9s�w��w�9����37?�X{n�?9>�͍������c���ɾohe'��ư��}7���JK��O�ݒ�G�%u(*�«��zo� ��hk)(���Dg�tﶇ�m�����L�]"����O}4������E�[A#�������g���߉���K��XO��<�v�vJd�\�O��ΝP�#Pr�`"q"�y.����W �p_:Ļ.T1�\pC��އHN�4�7�w5� �[���YoX@��!���
zwy�S�!8���� J��(��}��2KX��U��B����I��i%W"��I	Z%x��N-B�ؔBz�y�Y~���U�@ތ&����7���@�x�_J� t�zz�0^�C�mj"f����x�����^���p��)Ӛ��t���,���m�ZY7���>����2��c0�s*���mqO��?�Sx��O�[y�vzc���|6]y�<Ɔ��=3pG� ]���ŷ����w�����F�7Ǹ^�*m.�z>(O��8�{֭�?�B{�..���]��@��ߋ�G߈�}���`�n�3�����	Fv(�h���4>~?�1����x�����O"^xv�gt��X���t���w�?��}3�v\�z���f��z�D��GW�������L���?���X7s|�e�p�'��.˱=Y���y[p�S���Dߏ��zW._�O#d^�v5�:�25s��N~W�O|���������}�e7�C�*���������,���,��g?u%>���X�=����N�s�򥸲����������Hy��� 0����+|ВJvY���e	���LO�QC�cXYM�Ty�IeK�NI�c1=3�������,���䡯�Z��p��>0}���\s�M�۞V5t��n�$�pY�l~�mOkU���-T�h0:��ߔ؀%��A�����݊���>�՟���>���{��/�����s?Ó��Fȴ���f;�8���y,��[)O���6h<I�9�M��྿��Ffkd�L>��	���V;�k)��/��ʥ�[\�	�9CY�\�?����_y!��]Z��t�{��p*�$k�\A=��S(I���n��?�ʑ'�L����?�q�E��*���f-�Sl>�3Q�؅�%Pi"a��.�[�ޤ�erI���T�E���Ap�+<�4��|�����|A�/vZ�q����hw������4���I�D�W`�q���i0�u8i�ط.&4�5��H�״@J��#�|~* ]B�"���/�2�V��ޘ�J��d\E���R��3�b�{�wHvaL7�.��^�� >��O�5W�Y�/�G�n��?��ht���?���&��(�P'��X(����w�;��h �B��c]:nvQNiu��f�1vVW��Ӆ�Y�7�y%~�3���R��os
��>������~?Ώ߈Í����Wc��o�����ѣo���[q�� N�����O��G9o�	��]��rH5�k|��v����XZ���~����O2.�b}L��@i�$m'^�q�?��#��~�Xc|xK��N�b����s|�P'[q빙���lq���Λo���nLOv���|�w�m@�]l�M
��O��|��S�ݤ}�C��Y�VZ4�>��q���r�˸x�T����F���tyN[�L��l7>����?�q���p[�s��_�g��B	��Ғ�})��q �l�}���3����>�{i6A9�>��[���nѱ{�� 
4\i�'����ܭD��5b�=~x7~�1���/���~L�g��o�!|���� �jρ0�PpM��j+�Id�y�d2J�s@�|���)��2��*����q�.$��ܱ�՜��3��z).�݈���d\����=w+~��4n>�,�݊���1�ی�c̷��f��"M�/)��/��˦v�}zo�|u'��K�eG96�Z|�]�P�'�ל;�!�[�U\Qq�yc��.� f�gn��i�:MS�d:~���x--Єr_���2Y��X�n�mw�n�tk5�K_���?��A�Y�8�"k��.����XĚ���Щ�Rjq	�.�����L_�R0��=i)x�Ͼ���m�)�K�(�n�X�v�Kѽ>����>��U���銫���~�1�	@l���\o#<Ͻ��gӪ!�TZӳ1�p9��+њY��\�D�]���<��M,[��~��ь��([*��;H��~ev&^~�z|�C/�ҕ�1���G�����lO��P>D�|+N������[?���o��������^����_��^��X���J���cp�0��uHn�RR�=J�G0�c<+�#���&�m�J�*�S��X���˫s1�$ 1 �Ÿ���98>��Ǐ2�Ӏ-4�N6�o��J��z�9?�����V���Bf,�7�{����"Č't��j������L�9��3��8W7�������%	�*����=��2}V!ߟ�G��G�e⊡�gK>{�G~i����8���Oŏ�؏��囱�sۏc�ۊ�������=O�N���n�J�#r�����\.YI�o��O%(��.����1L��?��AX��ˉ\�?x9��⃱Hf�J���v�������o~5����3���o�LLN��R˵�i��!`,��k�"�ȕ�e:(}y+�4��VKH��/���I����V։����wNPIͭkD��z�j̯�`	ͤ���[��O~
��|�=���� ��h��d��;� O��T[cX�ʠ�V����=&�|O9ۘ�s�� v\��c����$~��i{��,QB���K��5k-�Y�
܆n?r)���'�tҤ�!N� ��� :IS�B�M�G�x�v��@�]ߞvgΘ�$2�'��{Z��Ψ�X�X�uP_n0����^���7}I�8�}\����:���|�8�ʺ�WřF��A�S�$��ɬۓcqem>���0nd�GА���iW�o5��H��b�6�Պ��
�=�HE��4M'&g/E��D��c8s�t�q5}��z*�&+�g^�[�f�u+y4:�X���K�8t��3V�MoV�l��5������(G<�l��p3�go�`�7b��_��_��x�K;~���N|��~1���8Y�^���V��b����Y��ݭ8�܌�Ǜ��ގ���������
#�l�yh�(~���w�ă'z��d�����?�Nq�}�@?E�l�����#��P ��]�*iG:Zf�H315�ޜ�篴�l��V���N���aU��l1�W�fPf�brf!�S��8Lx�.��13|{�8V%��j���dG����1�b�B&߫y����Eǉ�����L�_+6vd��G�Ў��N|������P /���.�Տ�K���%`��S�1Ĳ+�0z��G\s�8�r��T�U.O�(iJ"�e/�{�5@B�4Ն�X�����ٗ/g5�����_�����b��}�J�_�ʀX��yLt�'�棅�ќ�*A �O]1�dWss]ǝn�Ύ41EC��SN�U�K�BvJy`t��R�E�
R��q�i�.�����1m�=�޸ן��s�hW���&Pc� ��oA�Χ�L� ,��٫ΰNM��T PBf�y���Q|�1���6+R���Uٚ��3����!�����WU�O9�X&`��^���X\MXUX
�l0�"b
>�  �n�	�'�̀ә�T�N��$x�(�d?�cLg5>;�.�Us��� 2N��ʵ�����_OS���'E<)7����X��P�'�J:�G�,-���ź�S�s���;�N�e^��j��HMA�L�^����w�#��������16�\4�_�A�JZq���3��|�:�A���2��g)��5�b��`��l�fOm_@J�u�B�à���p�G���T�=�+�-��磝`��)�������~.���ߏͷ��XCk�`�t7vo��/z��b���q�����;������������7�n�l �:� |F[��xmx&��F�zR=��C����8><�{���>+iN��0l���~/޾�����_��1cX�c��qp	^J��z�|�xa!;cq��UZi�
L�֭�q���X���,.���jL�-���<h?]�Mwv.�y�
!���t�yo77^�����)�z�'?��F�@zx!�r����~N�c��g��w)�1?;� �d|��?g�N��,���ѕ)2P��"��zL���Z�x��X�Y�(._��_��}�����];�*��4�Q<	,��2(����������r
������������y<��V��>��܊��,L����A�'�q�b��d�@�MN����F ���l�\�*��Һ���:B=�V��PڋD�+�5$II��7^\��{� ���?~����@�����c4EG�;��QV
n�]ʽh��s�U�@����L����s��J)\����",-)w<w=��ok��uN:9�Z��9�	JZ����љ��%ȼy���e�Lz_~ ��O��Y`�D�Ģ���D��7�W��ۃ���dt��x��b?%.�G�dX�Z��:nDpZ��}A��[��+�����8u����̟�T�x[�]��|���d��'��8���D;��/�n�0/���iig"���O��q*�?E-e�Z�CM:���\bo��L6q�B��ñ�8o��t0��i`��S�[���C;6;����2;�1���~S�����KW�7�R=Yѹ�j��ю~o?�m�p&��տf�Z�G9jl�H�s�7������s��λ�M͌cx���<wq.�ڗ� ��~.�u�����������<&���_K;Fa+S��C���p.N�����r����{h&��R�ť�9��`c3����ͯ�V|��ߎG���3Z�-�I�~�FY���XL͏Ǉ>4z~*��G���A��(�U_�~%^|���~�V�-,��*�DZ��ML���^ޘ/R�
6��/���=�\#�r���xJU����:r�[�!�\U��ai:pL��K�vE�o�_5�b}};�ww�}���c�%t|'����\�$��p)O���$qJo֐4_"ݱ)9��D��eN�0���<�|�\��泷�^|��u bcg+���ټ�N�L-�ڵ�1��� pg�t��-d�z�}j��)��1���$�D��A�d�q �޷��)�H)3��)���/��y�T
2�$�b����g������u1�Xo\�Ͽ�0���m��y��!�g7A�������nΔ5��+�0������9a�%�yK��t����,��3�N��߉�G_A�ZL�܍�f�����r*�t�"�!�06����L�z,���+:lZ\�[FZpxw��b�8�܂�!��(�S��S����O�&�QVZcIk�]�s@nq����L�O����T�K"��ogYL�?<ا�t�?�����J˰j�UF�@AY����3ܕ	��*o��2��;���W�	ۧ��fұi��&�I���P��9��::D_%����)"}VT\f�GzMo;=�OfB9XJ��Gh�.�|���a0�G��8�`FBa��4�i|�ª=�f�`�|9ֿ�+��/��#�'i�&QR��ս3����c��bLμ����K�k�q�ʇ����`A|�>[ۇ����ظs'Ύv�a2ڋ�Ӄh�ֽ7t�v5E�I����~�������^��{(����w������ƻ���	֓8�v#�z��x�] ���~,�b�����Q��Z{����2��=y���byu5f�r<�����|}�[>� �j1N�}jf�:��������7������Ty�1��-=c�U|���l1n|9T�#_��b��.�E���W^������fb�S��嵙N,wFѝ�S�j�2=���Y?��Xt)�rF^��C��ˁ cTSV�K>�m;a~��s�W�ō
�x�w���z�m��ڕ�bai9�1��'�*X�{�<�h�8�EA<�$��0?�\��q�t����I"9%<r���VK�LPV���J�$n+ӳ Ga��v)V Oֽvy5~���b����N)@p�����'���e)�S1 �?�p5c,�����'��..K��-.���^V�0lx�P܎�����/���oFs����4�A�V�*yeQ��Q|ad�l��^(�H̪#��`�!�.w�9�,�G����&����Itm��4�kR�G'>H�b�}ƙ�8�,(��{�� .�]���J�V�WO;c�K�W�ml�����{���U��~K���@�AgU} ,�!��cթ<2���N�
��q��䜈�p<$Y׆�}�	[����,D���|��7�'����+�g�I�ő\P<mzss#���]���A�nh{�z� ���ݸ�;���[q�w�&M���^Fy�B�J��K��D�493��O��\�ϭ��^F �/�����v2���b����}�(�'�Ř� �������s�����,l*g=��[�{'���߈�o�Fl���;q��v�v��r�`�6�~.��Ps,�CB����\#&g���y ,�0쩸~�j\���Y��ל>�ϕ�=�V��U^�Ѥ���)p���k#���s(���+�5˜tͻ(���<g\�i|>;~r,��+�R��6E��������s�c��.�L�c��Z��Y��(pR�}΢��>�,ܱ,ɟ��>j�Y+�z����E�����rŒp�x��~|�7~%���V.���\��Y?��I�Qd�&mgJ�&Ñ��\���۴^�i9O=v�N�S>4�F�ETLK�Q���gb�8%��.&e6�:��ˤ��ՃȫD�.8- �:^���g��ť�O���-j��� `LF5D���׀���d@O�Igg&�/�	�Q:X���󒮤(�e���18�s�ޞ�����H���)�d3�{�����`��$�I���i�x͒��Qή����\�8)L-^� �'�'*��Q�z�e�݉�2m�}ha���S�?� ���Sj҅����Bl����*��=] P�<��?��N{�9љ�{O�V�_Y�NA��_)�I��TG~����˱)�+z��F�;����<N�s8<~S���(�$wX�n͙�j��#M�w��su�E�U}�����c&��r.�]5�짮��z<�8��BQ��9Ï��;���_����������vH7͐��)�fs2���j6g�����&��\\���/ĕ�/G����^�nm�����A���C \:8�Z�ٶ��6鎶���=�����Y�;�l��{�r˨1AK��||�|; '|��X[�O������1X��K��̳��*V���2�{���A�Xfu�e�嬍k�9�r�_?��k%��w�懥\c]b���v�O���
�]Ms�2#Q�ɯ/_�/��������b"���1�<��������I��Y�������!p�I���	��h�L�BGif�a5����|�FL#,�}�_���o��%܍g>��q�&��y̍��&���l�q#��r���SH��@zN�LwI�4�&�Bl6��H����<��_�TkP��ܨ�	���/ۘm��j�F�F�Ρ��,.����"0L���\|���u�n<؉88���Q��G���RB�Xw2xS+/0�{���aO`�Z1��}���AO�
�P�MdjZ�s+1�v3�g�E{b��l\���SM�'�����e��eWt�B������=:aK�Vg���&̙&�w��5�o��ko�!�-S1x�<�PU�-(��,E"�F��R�qⳖQҏB(C�`]����I�}������=VBřu;n��4��{$��h�&~+W�^�*�≺��|��g�'�Ԣ7��5�-=�!��B:�↎��<�#�mI�
�Ɏ��|kC�,g?�O/���r�c�����
��4�KnW������u�S�I�0��7��2�N;���xWguU:���#�h�eS\�b���b#�Xg"��V��s/���ba�<�w?v����n��Q��=?�q^Ɨ��G�\�����3���{`X9g(�g���8�3K��i�8���&�����鉸��.3�q���1N������7be�J��/EŹ���%��ﭕ���ėe��**ȵ�\f�R�Sleڮ�y���Y��ҧ���5G�uI��	�t��X��E��χ?��x��-�]�~yr<fZhz�"K
�/�����y L����N�GdD�5ڼΐ��D�S�|� �F`r�Ʒ���15w)��z>�.�H�,2�f� ���� SH���E*�S���4wǙ��yM߶͵!������Z����8}�]7��� � �_M�y���X�]�g�=� u�h���@���-�K�x��N��Ƒ��A�)Ep�\8�;���q�M�5QX�c�eiM�v���謾�7?K�..=����-0���b����/��b}�K�i�:�`~
�����vT�O!�Ʈ��R�n�Q��>�]��q�b��LaZp��_�.�َ�0eI����Y����eh�L��A^w���9�x�3�o\NePM�y���\��aٞ$0���U���T(�R�By���\��9�����)�<N���w�'�@Ჯ�SA�<�Ś�,�)�s����;�O���dy��6��i��XGG���o��T�Z�Ͼ��@����u�]E� ��X"�q�q�q�p3=���������9K���Z�/�NND��Z\��pF<�{/6����V~����$N���>��[��%q7����[6�ݘjc��Q�&��i�`�ܰ�Wi=�Y���HZ��t�a��6��c��z��Ε�K��|~���L����5ag�.��L�K)�����q#�k�9㣐A��R�$���<N�S��(���~.���q�Z�<�~�3k���/�d��[т����J��R#dl�H��\�Y���J��@2#��k��V(ٔ�>�/ݘ���p�4�G�����w�
��������u���*�]N�yV���NN�x��@p"� �����,�_:%?�L��^����c��;Ia�_���U������iZ#?��{�6|aa�g.������zm�{������s����Uh�L���(ڗT������i���D��IﴘL�n�f����G��_~!�W_���L�}�`��CxXd̮U��*.`Xz���&tV]��5|��f��#����(�I������\َ�§Z9A%Mip�f=^/�.�}��ˊ���R��(�pSG�}H�N�G&�M�Qcy-i�U�<(���)!b@��;Yna�X����u5��V�4���J5�D}���j���7뢻���E���3,��~*it��;`��˝�iK����\sr�Rc��8�~��z��>^��1�r%Z��c����y,�7wc���ؽ�~��~;��y#6�~-��'���x����i� ��Σ�f.=K(���~�l�ƣͽ����I��>��?�̝����D��� �N���x��ji���_��V���D�@�u*����-bAw��;q��C�=�vfs��,�o+A�v�����п�A�_�,��`|��M����w�9��vy��*�<՟��+��']M~�zl�c�i'�1\�w�ƕ���Z�]�a�L8�g�����v
��U���r�|
^~cH~B3���7�+����ˋ��?؉��x#��܎E�ޫϼ�˕@����ո0��^��MZ-N�)��ï���sԐ�A��"b�BH�*�=<7Ԛ�s���H��S���[�Rpd�}�q��t����G�zg�, ���S�<�T�ݕ��>�
[�y�3J��0���^�Ep=�qT%��_�=<Ekl���y'��:���6Q�i�
��H_�f��,��i��$�2�j��O���+3�������PA�{h�0'y�D����@q�&�`StPe%#%�	��	��	CU�����xq�g�1�_{�0A� �o^�\�1@� �]aM���>3�,uY�Ro+iJ�����n��o� �a��ˏ��$�ρ.�Y,9]w���z��wk<��P�x���ј���q+�)�87�򑣡Ж���ƹ�U����oG��<:k/G{�h�_�Ʌ���[����O0��z=ܾ���G%������8|�Zl���8���q�sRڠKNh��簒N4g�ĕg^�����ay��c=�2�r�%��t�E����ܾ��ގNsK�(��w|���{�����H `��͛(8���逯�D�N���|
�9~�./���BLϺ6�:g��������4�� Ty�;�K�xN��u��R1�o*pr�8�Fz�L��������~oz�gO;��[Y��4Aݹ�0N���p�)�:��ب�}rg��2�*�P��4<1^$�l��8�ܬ�j��Uj��W;�ßz�fm�a��Ay�~����ƍ�a1,�az��z��Bhx�9��b}  �����~�';��Se.4P��.�9�fz ��'�U7F�jgГ����Fy��3���Kt2�2�"�Ƿ�=n�݁�q�y����2���
�q2��X�B�f���x����N�23wdMj�j�fsCb��>�ވ,��>��z$
�H��2t|<z��.u���" ��O�3s�.�����'���9衤��>���0���OE�,�2����@".��,?�e?'���T�ܔ���wp��)���T:
�bh���;��4NvL:��p��[��e�5�U�M�^��N
6�������Ҹc��:Ri.��8r$�2̄��A���+�I�.�\����6!c��f�[X��S�<��.�n����﮲��u�D���S8�n~;ֿ����7~&�G�hϭ���ZL�+:(y��l����K�H�X�ƭ��ㅏ]��>�|<�bvq"�Oދ��ߌ���!v��8;�W�>�YY��������$��)�LL����^����"���ã}��0&��q����D�m#�%#8��s��E��n�[{b̏���~�A�X�-/.�B��$����e���jw�s	X��S�@�*^�����|�ǩ��/���_Ay�����Ogy§��^<g�P���B�\�=�����(fQ'�C�lX+,��{��,)��Ϲo�:�� )��	���t���+hB/^�B�)❷߉;＃��s�?��k�lπ��uQM�.Bbz���]4)��2U&�=Z�Oкf�T���a��F'Py�[�M�� �S �i�������}�\1��p<�aqy)�'��3�i��c��@-��LI�L&G��f�c5㪫a�����R�>��gH��*ʞ,���a�H��0G�`���\x�0T����������kgXo��H��`�$Ji�\e!V��ܻ��w�{9���-�1�v�;G�
7ȩ��ޅ�	����)��!�ͣeț��� gs���U�`F�A��IR�����A����8,>�ӋGǥI0�Z)�$��Jۥ�˫4G������ax��(ͥ,��A˳1��rĵ�8[��A����}��x�@~�9��p��g��8*x���q����7~=���ўʣd��NCq�e�O���/��f���������O�P������������?�ɸ���8=|?�X>�y}��Q1��v��/���R=HE��H����Һߩ�2=><�{�����D-ޯ��ˆ�����5�i>� ��8^K����ݝ�|�ə?��.4qy�}(���.��e	g���<��;������b~T.-&|�CXN�&��vg��?L��A{�c]��.]N�9����6�a:A�T�*zH�K�	��I��yj��ED�n 8�����X��8�Q���߻��j�Ώ�i,Dw��)��Sx�ʙ�+����X>�&���Ew7�@XKٲ���dLc'm���~.�qQ��W߻�7����w��nNyKZBd�� =J��h� W�zq_���`���^3��9���,���{��'c�]kE�7�$vtRDIsA���L��dm�2M�͹��õ�d+��2iM&�D،�����=�㣣���{�F]��̪?8K�Ź���# P��(4�U��㿂�0WcĦָ��*��{Լ�el����Ld|]����?����ařŸ��x�j���lY�ۓ�]��ՔZ����g��gi&FϯF��c�blf��v�բX����ߏ{w���G���yB�G񠜍���q��8�u�XT3�gU��s��D۩�r\�T{,�]����p\��O��'?ӯ<�K�E��W��G_�+���ڪۭ���ՠ���6�����F��z��*+�R*,�-Wwd���b�67��[h� �_���y�$�ʾ�K��W�_'����F�=�ۍ����󋻔� ��T�
��q��ܩ6=]xb
w��l
�s�Ya�:�
%y�)�����z$��ӗ�\���K�9<�����Ƌ������YH��0$�8�F7�P�=Jm�8�1W���N+�\��l}��(�3N7ŧ?�R�B�&�b�0�`]����)/�j���t�5�;ӹ٠>"<?�M�\[�}�z��Z �S������Χ�.1~ؗ��屼� |��X�PUJ�Ư�鐡��k\���F�O�
�{�d����*���/1y_��"?U��:��<�J��g)$��t�/\`C�u����YV���������$r���`C���<���2� ������� ������7� $�u�N 3�r����ce� P�1O�;g�
��N���J��KE���eq=;>a�;e��&�d�dz_���=ų��l@	IB0�Ge�uR�*צ}*)�?��#<�����㫴Y�\3�pU]��@�Q���Pųc��)q��5N��vww?>\��CO@p�k�B�cpz�e�I�?>���1��}�����G17=�s1~�Z��ǣ1�
����=W�Qj�[�X�q#&��BP^B ]�ؗ�
���G� |B�������i/g�ж�C<<ej���0�۾���D��It><�<Rd��*�@ �l`^���1O2��^/H01�R�'�-2񗴍7��_Z� dw����7������uO��/w'Z?��g���'ݞK&�++�����6�Z�/ˋN|U��\-�u�a�՝�hb���c��	B�˔17� ��uc��(>�ʳ��X<��Rv@�Q},P�Y����OG�	ajv>O�v3�{�ϓZ%L�]����{vD�Pβj�t�����52�.ZZ2�Ef��h�'�f0�`�3۠���p�/��D�x-u�	�m2�O|
'n%�RY��Qy3���>��sګD�/Wz�v��%AO`|��<-�pj>��*Hژ��̦��,�H�6�:��QZ��7�ERH�&�Y穿j�����n�N���\���
��?dWӃ0�9�Օ�Fg�������M�z�+�[�c�
�lG݀BE*
o;<��k�kU0;߿3=�em���5�x����`}җ��=��xx` ��)���ߦ9����8�a{:���5��S������=��O ���(Ϫ��a�R�;���9
�B��w�Kc�2=3�*�����=
8�x�^�?x-F������1v���ף��Gbؽ�VH��}�<�)�o����`u~N��K7
F�\U��.��  �WIDATL:��"��=�.�OҰ���X���T\��4�&�?)C��]k�͜R&��O�z�n�!R�,n̩�N�qF�l�FP��|~�'Gd�N���9��	-��}�s?Й���Y�?c
���W�C�m-�_5��J��	��'���	N"����d3�3�"x���3��ƍ5�`Y�)��}��yJ�4��n
��"zn~.�VWcny)���y?�xOB@�궣ÿ����G�e��}2�˽uiu�.���$��Zʂڰ1"|�Zg�e�	~��tv�֞�x��:rn�+@��7�=$d�F}�']>��l���<e7��������	���j�����7�m���i�ܖ*p��4��RԈ=��UeC�tN�M&��+�͝���܍>��*#eaUmZ�+�����<e�M���Zh��XJ���/����ݝ����'e
��?��s�S�S�Q�(��ġ˭������˾�F,'w�eY��!8�z�	� ��SI�d��ɫ�T!�Iv��:p��?ЎST����ޏx�^��{�=���"���̓��ʙ��� ����u�����#�Q�X����δ1�
-�	U�5��.�craZ ��w#�5� @��Jl~�k��K��~�g��7�}�/c�]�0�I{���&��?h�����q��Zb����QXТ|�D!�?�s����~��e+��^:�������سO��|�^ssFZ0x)Bc���R�Gt�:*�ܥ!vM���/3��@�9�%�L��m������<'�k����#����m�,������^���$�ba�|�4�
�k�$��grGTb��*
�I�K�k�d4��̶	���c]4s���.𵱈�����Ln�^\[�o��.-b�Ĵ�a)�<�x�|�^�����Y�y0�����(E�����ˉ`�s����.%a"X��l����R��ꁺ-O{]2�fA�YRf�\<�x_|y&��b�X�ܙ�J_[����7�W�u<��Ty��2y���p�C0@�l�t|��d.�Z���a<|��h���;Z�c=
9�&�ii#ЅWo��)t*�sN]�(�x�:t�.��j����,��fo��Ì������aD�fغ
�"�x�����VJ-�C{v2�ՙE!�0��.���	H/O‏�����x�֗m�Л=l�X�6s#��Ý�����v���NR���O�*
�����:x�yp'�+]<��[Ι�qx�<���i�9M�t��4�+
i��Q�(�������?��շ�w�����_;v׻16��h�^~q��c��7�+�B]�{|�G��i7�	t��-C�1E�t[���a�\��?����|y-��&&:;A��,ˢ?m)eY��)�pc���g*��f:Ց��%�R�]���Z�~}�cO��)f�4H\���O �zqG���\&�S^�{�*�vZ<M��'�5[��l��r��Qk=�(y%A6V�+��G�67d�s���88jƃ���9�r�n�v�T�����Q(4�˺k�[��Y���z�"�;�ܔ����������jA�O'��]����v��vAh2gE
m��_������qv\��&�*�T5s��^����j�^�J��~���d�.K��+U��l!�q�}\�[9}h��<]6�D^��h�~0��7h�@�G���soc7O���a�YoZ~�S[��@�A-Tt�O����qS_��tO��A�$�K��
݂.u����0T=A��S��c?v�s�L(�*��GZI������^f
޽z�'|���B6/��=Da�]F9�Y�3��@�@�N7�4��"[*"lZ�j�g��I4�#�i������^�q�^'4gg�8<:�����8���&�E�v��ڂ�H�hb�(�����JC�s�Xe�sw�iq1X6��������b�d-���h\��?�|&�S����T`,��9�8��x��í8>u����6�����_u�d[���a�s��3�9��[u��{{@�@$���2=��0����@�� �2M�L&#$� #� � �������\u�1�9�޹3w��~��9խDJ�;#�Z�"<<�=�=bŊ�,i�,���
FټPngF|�Kh��C�����)Y&��
�9Ȫ��_u�}M@-ipT�y4��i�@J��qα��L7r�
�[�&'����wb_�#b<Ugx9��}Dߩ����-�ɵy�N���oGfj?�k|ILF�7?��_� ƃQhO����O^ԏ?۬�S���-Dw��cO@��D��
K�Y*v?�y4���ꘘ�5��&��/���T`*�<����Ɛ�<��?:b0TqX΢�!I�D���5�-�|����ص������y`��J��y�C������(X%�6�ܭ-��1��@��9�cy$����9�8��[9���9JH�⢇S���ͽ�z�U�ݣx�*Y������x�A{"ն�!������/�Cq�/�����0��FՉ�kc���<��=�|�u�\�3z���7�h��ź�[�v� ��ƾ���������l��Ji��9�����LvO��Ey:̟�V�<���iGC�ۅ�'��$�)�g�W�u��g����0����imm�����ل3Ӷ�S�l��#�Ϻ cs�GA��fU6�F1��6�3D��rMݺU+������7�'���Y����U����׵����y�k������=�o����!��go볪�����;yF��b����iTK��.t���yu1m>���~����� \F�N���F�!����J��~&�e�4��*�Q���gL|���C�<Uls�r��˄N!<'4�Yѽ¹B�h��G\���o]�'41z�8�A�a�#ظ[��'d�F�1��|�O��h��O�0<>��������up���P)@�[�w8�w��K�eu���|×��.R�HCL:��
qtoeBz�iW��I�	yc|��ЈYL��K:�ǲ��<�|YN���f	�(4e8�?������Va�ͼ*��_����n��͔2�k����PN�I����,�Ɯe�Ës��|�\�x��}RKS�I�����S��$;2!8:8�����f	c�/��tD���z�;Fdo<�m����;(�S�ͭz��~��}K	:����z�A��vӐ�6nA��b��4��Ǹ�������eTY���:ګ�Ӄ����v��S �N�\��FaZ�x�TEɈ�W����t�[�^��V
e���?fc�ѓ˝��U;3��ڝ���N0�G5���;Z���S���agf�f��V����Է�����'����淫�ߨZ��A���F�%�/R�Ϟ��Q��th����`��͟���4>�:�1U��U��2t|��݉��ӌ�&kiv�.O����Y0r�12��T�'2�)�_��p�������v�m�}NII6U�a���1�s��;��� ���e�ۦ��A�)��5�ш�i�S�F�T9�fpl���fMP]�>��x�v�kpz�p�$�}����;���Y7�i��4!���n��g�Z0C�Z���×US�+���xv}<H���q�2��>��O9���(,��gi�+n��6~����2��&�-�<R6h6���&e���潱⍀�[)��=�s�h�R�Ql�{�u|=�G�N�@�du�����Y��h�Ǎ�,�!��Su�W���-<�u�Rpр0�1`W�8����
�z�����s�Kg����#�F�V!h�����`�Bx�G��E����Gw�փ�58F)��|�I'Z&<�'|�W�I��ti����k1� R^N�I���OjvpRsW��9���	�~x�Q	
#�+`/���Zn�A��W��G���$������v��˥�;�urr���a�r�qvt4�;I��jy�v�/~��;ݫt���N>�6�����E�A�2
��(4�ݙD�92��X���ɩ�<8/st:�3��C������|F�?Y�)�,� �S��j�Dƀ�g�躁��֝�u�u���Z\��M]����[y��L>-��)�i���;D����>n�]2RD\`����/r�$�h��D�������`[���f][��!�.���d�=d�^�5q����l�@�Yv�H����[�R���6���;xs�������|�,0�\\�]�O(�>� �)�^�ODy�f0���&6������No��G�^�j_���x��;OȈ��C�e+:�;����єySV�X�Ee�JSD-�`�WD{i؛�*��b�,ˌb:�i�σ���kh�=7��`n�$B�%������/�u�tLd���837Y+��^��ݓz�p��w��Y�F�:\P���.���<��>nSۺF�ӌ�x\��O8c�^�����i��.�M!����s:�e�O�=���/j�^�)�_��� ;�oo�5Z:+S�0��&����Y��q"ˮho4X���8MaX�Pz�x���˚�8��|�ɛ�c|2ϩ��1��#���G�.���!#Y�̳A�lm�g�;��ýz��Y=��y=����O���:n~��qN�~��z�֮���|�v-T����;٭�n#�e��h��U60r��s
.�#�C�C:n�s�!u����&)����?ط��y���õ|�FV���A�
�굫n�1pg�v���o�#�)D�����yX��63]3�VF��ȧ[�? ��,D���,��cg���Q�CZ�tNѽ����5��}�7���Y���:���צ�=3[��B�8�*�80a̫h;�V��$Yc���WY�QU�y8�(�S1�y��9\����Z����z��i�t�5B�H�8*z�m��2.�T�$(����c�s���j�������7Ut;ӕK�fȣ�jǃ��_k��%6�m�Xd�Frj�T]�?�#��1�GF%��Uޖ��bS*��w��76�b]���(�s"p<�6�G�(%����Ǚ�H���x@.�F1v.&��xAt=7s�Va�}xV>ڬG���J�����$��4�YqH�
�F_��\��"��t�}i����Fh�F�,G���{#��@�C G��R?ܩ�S���_h�l'O䧡j�䇣���(�lM�鿶\;�S�l#@�1�ϻ�u��B<����ZY\p��5�$�/a�6�9��L�@N���|m,�d1��Q{�s�������䣏껿��u��O��p8��V�5�O���Z��z��Fml���v���1h�>#�sh�w�Ct���Y�W��k�lc?}G��P�,�Q�0w�^_����i���Q�^��k��4α������Ő8]�m�Hwfía^��T�����St����٪~�8����H�N˷4�,����	��,"�Y�y���☟S�/�:��9Q�!|�`�BPN�\!WOܫ��5������ 1;���..p%#T�T+;�'�����<��A��#4��A�I`�=q���>������7_�V~��yLW���V�r��g�o��@����X���#�~��FD�B"4�����ދ�m3��k�5qC0 ~��-�ܐ�cE��IL�Ȯ���.y�$���Q9΃[~f�fcZ�$Gy��\����xzf����|Ml?ʌ�2(2	Ik7��QJ��ɒ;���Laxfp�g��(�r��m����j~�pqY�?߬�?~���!+{�m�����J̗M}�,��P.[�T�h#��i# �]}f{�|��7���8�`�쩻F��wS�8�p9�<��;�[w���.�r��e���H_
U��+0��z��8�ex�m�ǡ��"_a"-�_mj7ЦQ�s�u�,����o�*�#�9�έ(Q�T�NO���b�}�Z����~�z��k��w67�{��z�ţZ^���K4�_zP�� �r�&�Vk�Λu�?\�WutzD�s�a�����z¯��� �G���8�u�����YW&�|���[�T焛�0���_T-�]s7�W��)�d4�g��tj`O�I{�ؐ�ZYZ$}��m���vj���c��9e7k_������f����$.7y�NA�����ӧ����������:�g��_�?��==�����{�n�0Rt����|����3#�<G!�l�8���!u`:.�0�j�μ{^ $��QA�����<����lݸv�V��j�m�a��(?��ǐ|Y��z�#}���������D��]Pa���]=������ޚ�6���ԕ�#8��3~Y�N����A0�X�^��k����Hh:@�%^E*��΢�Z=��:��MQ���J9�&��RI#���%}�N�֔%*81����;�j�4>��p��vU�(�K,Pg�Xl;d�~x�>�k��٩K��/�˷�;��ʶ�q�����j��.`A35�CG��g���Q�bteBX�>�G�6�ѢC�p��׏?�[��b���}��py=��0�?B�0N�t>h��F��|��oyLYʷɍ�B�Jo��6��Q��n�pe����]!�,
ti��&h��-�>9߸/!{�9ewU7�'��;���W�ʗ~{��z��I=g���^_���k��MxG;�Z#(y�6ޝ�Z��F}���b��ƿ\�g�ux◀/묷S�;��h�a�����Sy�s2��<�/y*kF4���۩Π����a���W���|-��f�/^�9s�6���!^F��T�t����Nj��iw0]�N'j��qZ@���̗QזV��g�<���Kd7��b8�<�0l3�M	�����������`��ޣ���>� $4��>��^|��I����?�B���a�j�ؕ��o�"�5���F��n4]���H�!o_"Rʑ��pJmb���=��n�������r�,/1XZ��c��#;�A�AAORֽ�u�z�:�#t�x�ޗu�o��<�s��)Iʤ:�e^�~��K�3$D����U \yt��WO�=�}�	0��E�Twƅ6NE�,�b���-Tz@Kl�ʩ^�^�%Ͷ�0�\('T�۔��Iyaղ\�W1@���Nx��18�2\}��rw��B�OC\�ǯ�Ɍ1�C�QN�������W�A��h32���^
<�G���!a���d'�8G�Z��4rrQyև#�,�����o�w?R_|�I�o!����������Ԅ�Z��[�����*JGCm�Ͷ4��M"��%���q�ǭz���+�MQ�V.J�aé��Z������z���.��Y���.�0�G�PƺU`�q�����R�	��!�oA)p���p�r@�S^j��ܜY�By�u�jE�3')�Ac�����8��-i�2q�3"�LS�\���--�F�w?�W�ݺQ�|�=�����^�:�1pD�kb	۩f�#���������HMO��c�^<V*��#����U��E��6���.����!rL�p�cC��a��3t�]�܇J�����_�����ߢ�o���F�j��5�A�����^�'���u�w��C��1��Q��k�M�z�M�_���9GJn����>e�H��-��ܾ6=_��7kia9����V}��=F�O0�(��	F�M��$9�I���]����ߣ9G�ҟ��8�2QV��NÏ����Okc�~J{O0>�u��	�Q�SV���ZӼ�rI�2�H^H��Zg�ss�$�]V���>�;�G��Y��G�6VWjmuOwP�~3���A���%��D�����22�Z��V�������(�;��ﯣ|T:������ �_a�ίjow�v�61����0:�_��$�j	7G#�g�H������I�II;��s=�/�����=NWGy;���bɃ(̀/����@�����a����G�7)u�y2b2��4�3�s���{h�9e�|�;G�0��~������^�/�,����>���~����ѳ(�ˋ�h����5eC�����L;�.i!��-�w��BҸ�m��X����v��n��6w�?����N���k(�Wi1�c�h7�Yg���|�o��ؚȌ����د�`�g�!K��:}��^���b���8]�[3:D��-��		�G�2`8�κ�wt�czQ��A�|�	���曯�k��U%���8�̃�q�:}'_��Q`i�6�|��� u�~��x����O1n�K��V�Nv�{�����:�~P�۟�޳O�l�n]�?�֟��s�S��n�v��>������7��b�k�p�ݚ�x�ά0Y"·���$��t�o�E'^���IO-]�VK���5��Q�3�J�	��T̶�����C�A�r�w�
���mԽ�֓Ǐ���s�]���$X/�R:��ۨ��`5�N��	��9Ee��6�ީ������~��77���70���f��?X�#�(J�2�_|�sĄ���#�!���?Z�������ruZi�������q}��f=z���a�Rݸq������(�(�~ֺg�j�R�����aD��T"֐�`;ek�X�,��c�;����D\r�(�)�W�)�C3���<�0�rT(�s��i�֡k�����Z�\Aޖc��a4Ɏ�$��-P��їpiׯ����BtB;%mt�r�Zq��6��cGW�M�F�N�����/F�_Ѧ��)��Rl����zǴw$�^X���JX'����B�e�ͩ;�9�ڭ�Ǹ�|�Vf���Z��D�ׯ}��~���z��~M�zy.�\�|�]Y�O�$�H���ޤ��ƶd��6U,�[�L$�SZ@=�- �����Q�͋<�4��������spޫݓ������k�~Q����C�eϪ��. Q,�,���@î�-�F8r�i���N�%-���B/"��p
3�eρ��A����3� y����c�i?�V��U��|z0hϸ�$�}��D�i��Rݹ}����{�������7�S����	qT�+�ٻ��H��rfV^�;_��������_���ٓ���g����VuO��ctpquJY��3r/�p��겇A�>A�����˧������'L��?R��|=��g��4���F;N	�6tZv;P�i���e���1u�����Z��0�����,�%x7�p�s�]�@B�f�ip�����w�V���Z����y=�]Ϟ?��C�Fv��E�:e$�ct��W��9�������������96G�����/��z՝�^���O��`��}x�b�z�G�h:l�o#��vF@K���3��#��Z�F�	�6*����Ƀ�z�y���v��Sw�~��I}��'u�\FeC=�Q�x���OQ���eb|T*Q
�=�GS|�ߠb'p�}?�K9Qo8ߘ�� ++�D�_ �{��ic�t��[/�=��-����֎{Z�-�E�2�D��!}��,�����Nn�(4&��W-鍖
��c�i�.�Z"��H�J�L�F�
�Ϻ:=���������=�*}�˘6*����Rw$��	�<�v_>��B���sG>S8.x�.Ͽ�NԞ���]�jmc�����\ԋ����~Q����ųG5ٽ����lZ��Ԣ\���)���.nɪ8��Q#4n����B0���cX��{�=*C��y��:T�~���2=�>;;�'/�����W�>ܭ�_��_g$8���SR�������lqT�;�H����W�ڣ��ԅΠ���^<��J��؟���H�wR7�,�i��x�-�k.!ל��ͅ�y����яT/�7k~q㳈�Y���q��}�f���Z`�P����T�8� FJ��g_K�0^�w��g����n��?��;����h߯.��F���_ܙ��.,Pv�8�����������7j��?Z���3�q��Z\ZE/��~���qϮ���R�L�-�PԏTN-���u��S��?���U�[�t�%�յ�|�k����,�7���zf�k?Q�1��u�-�Y^���%�6Y϶v�����������fq�8��p);����b��1�Y�3mJ@�ýb�xX���>}�n߹��_�΁��8:��鳮,u����,���4$L������SF&��oݭ��c��s�"���x>~[ߩ6?%p�0|m}��ױvt��	���++��w�R�72�o��;����s��D�f�F��~0��;g��67	��_6 cc5㸁��
�ʎJq��w����7�!�����z�l�o`pn���P*H��j�;`��)�H"�������cc<1��B�<鍑�_�p�L���q�-^���p�I����r_�G�$�=�<Զ���ʈbj]&D�s�~�z4��rN��E�p���B�]���]�:l���fj~~����{t��3�)u�g�����6	 ��C{��6��8O�����X4��I.^��-y4,/Uo�*�a�j��\���~�ӏ(������}^=|P���G����{L�W櫳��G/���t0��$%���q1^9g=[�U�涵�r�Q�i��֨Tp�I2���|�2qq�R`ZG{&����j�=�|V3U��������on��ӧ���}�67_d��k�<�T���4_�~�m��4<m��͎u`�I��t��E6]�v����J����,�DǬ�.���]'w�;���	Y��ӧ���?�O~����GO��΍�\��u㽟��o��6[d��Hsz�Fsjv*# ��OOΡ���{��i}���k�$srv);���1Ns��8��y���g0�Ж>e�_1`�)}��qȑ���I�U9YG޸�Z� Ǖ�e�s��,#w�W�59�-aN;�a�:>��pPfZW�_H ������������\�������-�������,��	v=h����<i�Q�|yA��O��?�����I�g��Iu��xw
��c�����E���C���^7ո�n�9޷�ZYY���n5�M{_áOւ�à���);���Q���I����1ʑ��ɉ�*��+a�dG�GUp���x������Џ�����_G�������O��y،5�｣�Q q�g5�/�g��jI��M�Uk�(���eC�F���S��������EM�?��!��<P6�tĉ�y���ۙ�~NݼT>-ZǗ�Ɇ�H:��������Ԓ=���TG�*T��Z���i���;�>b��w��Kʗ��l�19z��|��|�-����aҎ����Y�^���^��q�{�/���e�=�{���� �"�/�{uv|P�7�գgO�/��t��}p�����V8'��qb����+���j�쵩����ۤE�s>��gg����/G+�����J�'�n- �e4vq�Q����� /bTn��Ps'��ѽz��Q��Y9���Z�_C1_e��)��;`�H_�ȴY���W�����%�m�Ϩ�<��u�ƍ7ke�V�L�����|�a�x��v_����A=}�[t���z��Y��z�;�z���?X7�ܪ���ZbD�)��Ʊ�3�3?�6��qQ��t����|��'�K��/c8�p��̪]g�7����zz�WG�װ��z�}R�=�������-#��mU�P����3ڋ��]������X� �@7�CGw�il�ys�d�a����Q�?�����Ud?i}E�qt�[�o�����?�Ӛ��x�f�pN���y��'dRf|���j�!��"�6M9@C��������Ͽ88���+��~ v;��p���C*��k�����|]_RІ��$tNV�������J�k��q'uv�͜2�!"-��!��#�/�O;�	�jQo�wDd��ۦ�����x��5��� ��rO ���'�w�W�.�y|vX��{V���0>�|
Ovaƣ�ZA�[?���P��F8�:��88�����?��MZ�����{U:�d	7�
���A�}�Vݽ�����v��bg�V�N�Rܦ��g,������cN�Y�=�|�c��X������9��Q܎������Ņ�ZP9�ܶ�;����GG�Y�:?7�QN�f�#�Ǭ�G.8�f>���w�D��v�#��̿&�^y�U�^w�k�Q'c8���3>�ۭGϟ����곧[�k���ߩ���ե�,��ax�l\���.�	z��k���՘a�'�!3�(F���Y)c�	�\�A�������;B��Di�x�B�3��q�!��׿�ӓ�:<ة{��������:8Tw8S��N=�;���vb(�߫�e��"�fҩ�n���g�EN�)n���0=uU�K뵴r��B��3"�;u���ɽ����z��a=���v��p�|����c���ڻ���Q�ɹ�Yd�����P���d�!m��(z�y{�i��_������?���;��|�������^}v�I=�ڭ�Ã��{�u\6O����X��0FJpϥ���Y��y9��\d)�+k�u��kԷ�w� }xH�>N�.��ᓽ��J��q��=c�ʞ2c����/�}�������z}��G����D�o���D=����yW��{�$Q���czI+�2�t�ɟ����Ͽ�?���k���#2f�4 ���h@�i7X��٠[�����Wgc��'����%����<!�aN��DV���9�H]ґm�^Z�����ИN����Ț����1-�&�e�v4����Gl
vXO�<���7�~�Wkw{�^<�gϩz�+(����R�x6��u9�0���B�
��a���4��^�ݳ���8O.�'��Si"��-�[�����):@���7���//����ƍ�Z\�.�
H_Σ	
IF��$6zr�&+1�d���Tf�g����US82�@�^:���i!1��q��x01��)=�Y���b�'�:�s?;<�����ǈ:M�🪉���n	ڈ�4�FV�����ܘ���G)��v�_���M7��� ��q�.·�����>x�>{�>�S?��U�cԳ��~�7��1<�+������� d7CVim�Y�%yT8�Y�Q�#^�,OԨ���d��K��OXa���:yi�UĦ��0z��ps�j#��H�x|ح'�w�����I��Pރz���d��~|�����v}���k{�n\����}�u�WW����r���Ƈ��ƿ#���}H��㲿U/��Z=�1#�O����_G[�z���2�j��T��?T_�ַ���mWx'%�qJ a�B�G��a��N1~5����f�������b=qT;;�u��U}��_w�֓����?9�{������zvЩ�F=N����)�����Z��o���It�t�Q�=�����(�Y�z>C�0����Sd��~3�|tQ�ì�O���y g�v����`~�a�'��������{������L.ճ��z�ȧw0O�рnG4��fТ��yG�=CM$F5�\�)&��}0�����q���b,\���Ǒ+���ٱ�:JG�S�����E��/��f9a�-ȩdii)�3繏W��_/��BH�=�3#�z�xy�|��ع�<U>v&���i_H}�PZ��>^�&ѡT2b���B��CP9;�ؼ��_���u�޽���F�l���;���˥�<�[�u�h/J3��/���	������7�-6c\���h!툁e~�Y&�@�2�v-~���/�^M#s�*�V�Kxsxi�6��g�l�����]��"���~�%����*2�b�c�wX3*�*�Ψ���I�r�
y����vmz�������/�+N��	^����,�tSF7/t8?��w)���j�7zJ��H��w����8KQ�##��'�1�7�kʊ�����;����?�>��>g�so��>x~T?�|�^<:�I[���
��ޱ�ߴ�Uڜ%�����:֑�A~� p� �D�ٮm_;�!�<F�gH�K�q��(m�l<Cɇ�@{�� �%�k�x�>פ�dON�s�Ӷ]�
����З�}��{>S�Wsuz9S�/l2::|��a��ռr���k������~�?~^�=#m�6����g���Hjo����`�y��lC�_��q�S't�cWk#�kow�w]T����/�}�
������`���zt�����׽OT���O?�{�����o��?�����/2�ڇ��57�d�XG���uj�^瓜Oa�1
��M�r{�x����H��3:��Ya���!͹��:���-���/u���Z���tA�%�e�(�~��o�VY[�K�����92�~(�|>ε������lY���[l���6Ev�bz�����������ÿ���K�O|�v�n���p�6{�{��#�lkS@�G%�{���h�����е���~���������/K��c�pa��(T�t��.?��o�Կ��������:9:ȧ�s�u�����w~���?Y�نg���N�U��Y��=�1��\�_�U��fܬn:�%�v.��2s�;����O7"�n��4DnLj���i���|��ѩ�?�q��?�����׳�볏?�G�ķi�1�v{��^���۫�tu�N�U�zl��r	*.�Ff�?Cэ��8�7m�_�Ay�c<"���%o�A��X�yЏ��J���:�Bi�o�av$KQ��K��j��:W����H3��Q�J(��� ��x�H	NC 켨��p~ʐ��������c}eXo���������^m>=��ޭ��C ��;��|����7ޮ�o߮�k7��Ud�Q^��8)���ȡ�lqe�<�i~n�d:��a�Jݶ����vIk�Tn�2����W���Y����g������ѣ:�K�����/��I?��114��qP�1���4�s�C�����w>�0�m�ӡ_�9Q���L���\r\�-�N�'�Հ:ig]g��ծ�x.<�aXV��@F]~ƚ3�ι2#\��K��[�y�YW'���<��^��r�d����,P�q��T�S���bX7p~�{�Z����������8aa�V���N��ƍz��;u�u�NW���0�Qm}zP{O;�Q�
�4��5���ZX�Y���ｸ�}&Ϛ��C����7�����:�_�;���A�Kt��Q�����8؝w�r�������\5C��m����I�g��Y�!+��΄������ˈ�,� ��Ս���A޳g�?|�{���?��?Q�_�������w���Y�A�.<��;~�Ar���,����|�4��Mͤ)�#=.$���O��}� |��iɡ�x#WX�s�f��>������������>��i}�+���7�V'�X�7���z]� ��|�'��i0�[Md|%�ъ�Y��|�s���������/~��:�s����h�E����ts02r�$���kmu��i�ۄL"�*��=����K��yw�����IAĒy���]G�;<��%	horj���q��p��v8��Č�J���~D�v������x9��zt����[�~t/t�P2[u6��t�N�0]_�ɛ(>�[>E�=�x;q�8��o�S~-�q�W�;B�Q7���-�h��Sc�mi�fȅ����6��[s���ُ��40IS�Y��9��4իi��k�%i��e��KAz���ʒ���~�thxy���;�(<7�X_��h�v�T�#?>8?A����_�0
=���c�E;y�Q�,�&�dJ�(.�T���5:K/p��YA���$'�ܟ�k��1<�?}R�~�Y}��'yޱ����_֧�g��������ibE���>�Ҳ�����϶��`�pc�yގΓ��(��4<NEj||��6��6h��|ӗ�u�|�6������$���|C~X�Q�I�sv:C�Y"N� �4���1~um�T�5���� w�տ8����z���>\��������cFHg��߫����_�V�~�+��[���������ϔ�
N�5�1��;�rg��s���~�^����:ܬ����ڭ7�7o�W��Z�~�upzQ����::<��݃#FaG�:>����ܯ�p����ۻX�i�Ȍ�~u0�5�O-��0�?�q�mE;GY�4�7a��:h=�����w��í:�u��!��J�-�f�ͯ;g�Q)?�PuiV�ٝ���@�7e$�?2����-��3D�s���vt��=!i��1���W��~��o�_=����z'�
�o��R��V�{�9g��)[�>�e<�6�V`�3J��5�E�<������3����:�S[�����"������%�����˺���&q&�Nc����u�(��S\�-t����u�K눂�y��N�P�K��wy|��yu(�l��g����6�yT4�76:-�#yT6A��ұ۹�����������?���������>]�U�T�l�:s�_���Ύ�%U��A�Z�s�C���v0��5��� ��y��"@[[^q��W2��m��DM���`�T������,}��8������{���kC\��Q�T���iĬ8�2��r"T�o�;���Co�������XOpn�i~vay����4��S���;����Y=�ޯg��x�[u|�(jpF�tQ�Π\}^���<�,�v�M;Gm�=�BW���Jڵ5n��==����z��i�����{?�a}z�A�o��l!����E�����
Jj�Ji�x�?�-Ɵ�,o����Dʄ����'q�z^�3[��ޗR���1Vf�\�}�%X��[Y����L��S��-��r�e.����R�eTO{&�1�s����җHGa�*i�T�(@@�h�#��e��!�b�(����u*P��0��f������{o�^�u'ψ� @�1v�׻����\1�]�U���׬��-\� \���[��9.�Yk��]7޺Vo��y�Z�y��ڸ�Z���K��Q��B�������p`�E�ި�u��Й_d(݃~O�\H�gW�����ʻ[s5��$��	���^�;>W��(d<�l�`�,���l{��|�{p�v�vq"α�ӵ�����*P���j�����ɻ8~S�]��5=[Kњ<�#�#����/K�8:�@hr�UKi��*���'�������[�o���[���u��ƍ�ڸ�ZS�uԟ�G�ep�9��ب��OccT�K�k���F�Z:A���g��+>��c�MG��َ�Ҹ����f�
�A��Cb��0Q3x�����9=����c����wM���3�AT�١�n��p#?���	��y�ޗT1@~eԇ�!��^nT4��K���̣�gY����_��?��{�t�!����ޤm�tN:�M:ڭŚȨ�Ec��j�.���qh5������6����iٽ��о�蠑��/5��� �.����[�$a�ڴ�rzSXN���r�g��R���M@_�q}�}���$�������L�6��S=fr��8"@�\�zN{�}��s���^Zx�~d�>�<v����Ç/�Ǜ�l�E�@7��0T��Y���=�����z�Z���3��~,���������b�������������a}p�~=�!;�j�lXOϪ>:���[����7P0�������iD������uz�i?���.jQn���D}H;	G� ��Hб0]�ƾ�;WmǊ�=�Ւ��_xD���w����8��dnv�i�vC�ǎ��0(h�})t��Rw������B5��_͹y)�Yo?�5�NK��Z�Q�c�{��j��y���Zj�t�-gɽ��8�ܭMo<zP�}t�~����޽���A}�7[w�g����z���ߝ��\�ߜ��{�zv|Y�\����A8�A9��67�W>~\[�T��1�o����5\���6p�Q�Q�hԒ>��8�[��`|�YFc�
-�8�y�o�{��1� ��u@7dJ��cD�FL������v
�[G8䏞m���>N��Cl�/�;]<}&��)��F���s_L�u2�87=��|�CW"~�@#��G��DC�˦F�@����֧X��K��~���~�׾_����on,��UF�s�xV��L]��Q��g������RE���GN<�	9Wf�VY�e�tp��Ϸ����b�|�K�B}��I�&2!�s�������Y�&z���-^՟�3_�ҷ��6N���|��쬇u�oܪ��{�^�}��6^����p�K�]	xr��
�o ���m
A�f�a��Kn2j���p�r�"$z��3腫p':���͆�w?��~�{�'�_��;�z���_ޮ�S:

���g�^��e:�Qi��sȍ�M�Bj.���gh���L��h!M���Ng:"q��(q��Y�PW�;��j�
	�TϽTV2Z4��9���ΪIi��v�h5U���Yr�(-[�&H�2��8���������]�yQ�P�u~P��	�����id浥�z}m��Vfj��?F�h��v��X��A�NwP�W5=�R�7���ٺ�:[�6���k7�ε�use��V�HW���eչ����У��t�R�����ۯ�]��I��	N�;
L�9����^��_`����1�n#b�qZjE{�\����^ɬ��(�i��+�z��9�ـ�NR�f��oY�o2ڔ�8�����e�m����������\���-O�Һ���#�%y/�O�x���L���I�֬���J�T/Q4�j�>f�Q�|�/�������(᜾r�t�?'ݓ:��6MLB��%ڄ�Z���7�@S��A �f�N���NN^�EC7dl?��.����K|bٮ|���}�)�h�޶!�u�~�_;�~�1���9&ګ�;{ �&�I��/����&�wǏ�����1��!��nem��ܘ�����=��k�[Z�^o��f}�'�V?���]?�s?Sw^������DV!�i�g�M�1D��mϑ����(,����j�4d�႒�]���%�3�u4u����֯���o�����f����_y{#+���^�>=�����MIx�]R_N+�p��e?��47t��z�i��.������7�n֟�K�v?݃� \a2��-�ZP�>� �Lz�Te��^��O՟|g�~�����Ԡ�`�����0D
�q��{_�FݺuϤ���*��<���t���L�I2��>�Y�j�9���@5�T��׳˶K�۴YemP�|n���}��I=zx�>�����/�@yg�y}�t��nT�s�w���bx:>�Z�p}V <��`)�(���m�PD͓���$O�~�QHooB�	W�IE�4_M�4��,�Y��J����CZ���#
�x���ֶw�8yU'���'I㩫�g�3�cg���N��.���Ԕ���w�MGd(1?G��M�^���4S7����A�.��uzܯ��n��2RA����:�V�,�-�Sumv����:��&+�˵���w�u8�q%���1���{Q=eE�7;C�Y���U���.���}t�	�/*_Z��O\[h4�b]bT0�2��I;��}3J@���f�����>�t�ĥ�.)O��D��EB�Iҕ	�R�Ku����.Op���ם����4[�}�N'��騎adX�K۝��S Q\(�y�ݷ�-�.0�&��9b�3SH������iG��s|/�"�F��{�u�{%Ȑ����N�����t����GWW�0&OP&�5�s{�b�����b�fn�^��U���S=��n͠ 3q��nӁ^�].Z5 �D�9����Y�~�H�n�P�؇�9�G{b I�鎸;=��#"2���D#�<������3�<�SW�0B;�ƨy~%��}g�~�g���������y�6Fk#<��]F��˷���G>B;�8�3Gt��g���R���\��^u�s���O�l�x^�|�I=x�>������6N�dm�/�=���:��z���9��i�Q0t����¯u��FC<T�3~�龃�&��*��Ƨ����F>���]۟@:a�Xd��S$znx�)� �p�4X����]N���D�O޽��yGa_�����xP�)��olԛo�^�X���u<�E���wk�{@>P�J�7��C֌�h4@5@���j݇i���+��*�\���Na��*�'��Z��E��٬��^�������h�N�6��O�xW����C��I�@<�([~P�	�J�z��m����b(a�L�.c��C��HP�e贤 �"�@��K]L���Ұ�R��'+Fٙ�a~��c\�����J�����G M����h����TՖD�f�4i�,B���a�%�_�x�u�P�wH&_^�1��� M-N��R���oq�>���n����8����4�e��Sw�u��&�0�v��r�㋇ˋ�P**x;�`���0?����r��Y�m��
�8����!���v��&��ϲ��ϧ�@�.��L��'���V���w�2��у���,���g�U$����_јseg<�o�#]�e�$�-���|g	�N_�j�|����8j(	�쀑��v�3���o�ߡ�\5=;Qss�5O��Mg`Ӂ~ӌ$�i߯�����[��%�y��;�wU�D��2%�O�t>B�|���;s����+�P�*/Gr\PY�>n)5|���N�>m�M�7k�οP�o�d�O�}|-�A�����X��]d�'xj���2���t7;ltp,�8����x������@jHeM�@��X1�~���C*9�P2j����}��6U7ׇ�v�_��������hpe}����w�g�[��o}�����ѿ�[b�8���z'�����>'>�6���p�_�]��/������䨶�<�/���}Q~�q�����"�n����t��:��_��ԧ�K����Wp�FG���C[�>�y+=�g҉��F/ŝ���5y�rU���������Bm݇y�T�sg�(E�����l�ҲO(Xt��3^6J���e�k_Y�o���rx�Ȁ����K�߸�QkX׵�Z�~���(?�P3�G�\�q�W)�"�*�9dΩ��p7�Fs�Z���p��K�!��cx�?٬��=��}������������ڧ3ux��m5�R(�7Wkr!�+	�˒];� G�Q��r����ު��(�_��v��2��YĦR�(6��T��Q��}��l]�S+��*,�oԴ�E^nC�gi/�P�(�H�S3�A�M�!I�t:�p�r�һϳ,:�G]yr�GB�|�'�(ȗO�����vi:�氆z�t�s:�#�����#�s=r�s�ԃ,�C�4̠��
׎���kz\1&TV=:Cy��y}r�'�Q}G$D�����,}y��C3����lw��ecE�ڬ�t&��@�c|\��7�9JK�z_"S���Ay>��<#zH~*���	N�a�J�Ws}�ֳ�|G���..���u��l���p1D��QʉFq��VS�9`�yt����-��:N"m�=룘lH�]�#)�W6��i8a�;*s��"@q�l,�jo����8��ƏW��*h�61yPW[[u���32��s���[����Q�]2�0���Н�B�B�g&n�{Nlȃ��QM����N�֮����.�U#�7z|�0_�.��gsE��e{X��#��"D~����3��_Ne`�>Y��:�:�[�}h|\{[���,c���Wߨ���f���[��o׻�}�n�����d�[��n�Ȑ�2�I��E߻�_����F�����������u�������'ϑ�A}��ku���<�� 6����d�����S�;#M����8���hVS���3ψm�4j���Un��vt��~������o��#,�O{c|( �4>ΉfN��
�t�Sv>�O8,C�߸3]�ҍ���k�Z\ҋ2��{�����ϐ�"�y���Vkaq���°�Ό�11�B�����֨Q�Av�fo[� ����o,-�2���{x��i|�������z�'{u���?�ԃ�y��+5ܟǓE�H�7�l�2,f�����@fc�i}��%q=��f,�u�=±��l�Qn	d�0%=瞴��t��y`�ʻ�g�oy�O�OU5������++�2�	����d,b��m�U�c�7�8�M����9���o�X��^KLO�؏��{C�ɉ>^'e}n��gy��+�� �c@��:Y7���CYN��\�L���_�:�(��u��#�'��!pxQ�'xs��-?~ǈJp�����#����#>��5tTN!��ЀN�j�p
1��������Q�ұq�j��̌h��xaJ�=s���iQaF�����6�q
ٟvW��-�1�Ah�t�f]�ެ��K��@c���EP�}6�W=3=�R��5���;K����
F�6N���ilF������/+�B�h�>������6�����Rm�ON���H<�ho�^����V䥷U�[�T<�ٵ�u�'�huު���(xq�U�M�
8�(�-8�S 7;ň�v^�����V-]��F�U�)�����lbgCH>!򞔽��6:�"	\c`;��r�<u-�ǭ�4�3>F�vQ70��]^�1��:��y/F���m\�V���Z��ʍ��;���i��y��yt'#z�{[^Z�jG�����_�e��W�?xVϞ�`ĳW�}�I�������u��O�,2����|���ȹM\O@����zt<U�#��d��@��L�ii�4��xu�	i:d�n|=��7�P�����ώ��d�����юX<Z����] �W� D�&,;-e�g����u���ʰ����wo�׭U_���Y�N�,�8�p������Y�����5��R��+�~C��~�K��ܦ��"�N�̒����)7߭�1��^ghC�ɳ�a���}P;�[�9<�ͣ��w4]���5<D���j�o��\[��9��]�ot��j���9�s(o�����O<s��yo/�N��q̦�c>���3���r���d6i���3�'�˿���%o+o�D��v�7x��;�l��qDt>��A:*Č#8*���	�Q���TR��MC����Ƃުpk����{�L�,9�z6-�O3@��ј��yF�t"G6�N������^�1*`��3yW�w^8L{(՝�y��%]L�U��8 �(B� _��S�}�,��g\v�4��"��J��͟�@%�T�(-���lxEsx��zl����Ѩg�fg�~�������)���=p�����w}�� O���F����{��6Z��ڀ�z��3(g?%`�w�G��"�A�]}p��ucF��gG�&i|�4et�gt�2�JF����,� �=1�~#�{�����J�Z���f�w���i.Y�Q�ѸP��U�6�  �L�.}�6{qTS]���zn��6��`f��Αh�;Z=g�O������[���s��+eN0085>�r����&���?�kk�um�W��Mԭ:;�{T�~'�fWV���Q���ʊ��x��WV��G����Ν[�>>9܅��vN����1�yp�n}��O���'uF[��2mx��;�FX�3��Y���g�W���d=�j�)��(X��M�h<�1��-�gl��5<�.��#s�9��}	ǩsr|z������Q[�O�zdj�
�Cd�L�Cf�ޞS����S&��x�֬��Z��ϽvU߾өחŠT���n�0>��Z[[�k7�Ś����e�L�!���r���fX�T��,���[�.F8�߫ϟ���v�h������{����S�g�uܟ���T=?^�)D��:$���x^_�v�>t�ڙΓ�4�)���ha|nC~�	l��Mhג�v���D99R�bj E�ĖE���*�Q�T�Y�ڂ��9��%Cڸ�v�i�DLy��?%^�&\ɝc�H�G�~;*�_͵HE��!�}V��wFB���ó�^���"�����L��s�N��ygi���<�2m?ULG�D���.u�.�j��*V�kL���UY���7[}w��Bn�$P@Sȵ�!S�$��������8��"Fnf�ϗh�U���.$� �,�iBC>���LGGy^G1��֞A�PȾ��� u�sn�/�n?���3�KF
f�����O|P� 6]�g<�65�Ne��9}v�'5)Q�<��I��k+n��������u@h 46(.�ZdQ�P~�q8*Ѿ�^�D��a����(���gh���O���G���ĀO[�d����.OHG��pD疣��}������J�+���V�Ob,?������|��#v�����͵v�uv�ͪ�7V.ku���0T.R�h\pt���%����#��Q]���ޛe�����o|�������z�����X}�����}�k?x��>�E$Njf��|��Z��Qo��Z����ݥ��T�߽��'��?��6��ӯv���Y���sT8"���9�j�Z�D3��^�k ̣���>:�?����قXx��x�f�{��YI�y�ra��U�N�0�\��©�_���(��ݜ�oݺ���N8B�3�j�gg0 ����k�����*[��=S����\����ɂ��w����\�|#67��N��g�`�	u�0rP=���g�6�����\����=�����LXsݾʒ�K�9�s!;�/���k$r�7�Qؗ�t� j��q.�M���w,�H7_�x�1�k�����0�-//r�~����.���85Zc� ~-��p���c��B��n�?�����G�ً�k�N�L��nɴ�"2*	�o�)c�������l� C��ʢ3�EN�0��ܳH�܈�j�R�)C�����6�g��PhT������!]�<���C-�+r�ma�8��"�S2�t"����*$��	,�G�d$�M�Shc����+�%����f�Qh�b�����T��4���@
<��,F�~�/���O?Y5�y\#C�k�P}����i���T�\\�v	=���j��<����6u΅��G�'��G.P�;�",�e�V�F�����A�%͉���E1�Oߺ,'\�P՘f��p�c��8M��I������	�-�ܥˉ�5��H�;�-	�Ӻm��֦�L��
FNU��Ro�X�o~����d�|�N���Y�͍�Z�;ǟ:b$��~��ZF<�g؛Dϝ2b��N�Ha2/�^m��}���Z���~	���_�ֶ�[��V0����o�So����_Ǚ_��3ux>Y{݉z|0S�N���q��$8ٻ���y�C��՚)���D��=F�2 G���HwE��`��~��^����7j{��N�)0s���6��q�IT�`f���|-�����}��� I�꣙	��E}��\}��D�MØ���Y�XoG/��+Y&�4����.����!�i��AArS>7,�A���~a`�D���n���Ì�����@����l��`�!��y�戇�F;����r%�+��:��E�]h����?�@���C渣��%�4)���ݔ�M��H�Qy������ȝK�-C�,��7E
���r�5�|f�6��P�$��3�sަ�,`�y,�5U�;�Z��o2]d>z�N�>��~m����%.�Q=�vE���yF�::��+:D�Ky�f:�-!�'M����*�h�q��C��F�z�������EļN9��}(o�A�8p?�(Xxi�D�0ãu��8XG��x+�^]C�$q�ғ'*T���5
���/���Ai��W��oV��l@=/�"�[x�U�T(�t�q,�6B��)܋\��eK��9�UE�|�:����G�tX�D��ܫ��O��q�x©R�:�@_EQ��.�`utN4i�M:úe�
�:l���x���kEK�=0�� P��A�����ᘼ�=�G�ς��ض�:�����d��7�ɳ�����Ꞑy��sU�D�Ϟ���I�-�����)��G��~S0uP�fQ��
\WV�kim�v������V�N�~ݹ�nͮ���z+�P? 8�������9<�����zĠ�֦�1�y�in������[��(ql��$m4z>�c����}<�#a�[��999��u�Ͽ��j���R�kq�h�5*x%~{q�^�.��CI�Q���aA��=ܭs���`�Pч�g�
�=�ūZ\��{+W�ε�������dm,N���8G1�e�ב�kX��N�w"�VYE�����EU�E)���|��63�v܄�m]��&"�?�����ju��W�r��(�yb��'�؊���+�z�\#�}�r��(���k��ܒ�怙��;jx�9h�'�+��O�7��DȹM@"���c���ʌ��o���n�������
��/A�a@�54>1*�4󏊤,�s)n*���Oa�㷇Ϥ3:��a����Ί/�
#�����
>J�e�0 xy�q��9�v�3:O਷J=F��+���{1Q>Q�
=o��MI�X.Q�ំF��m3�����$��͖�VϘ�-�nZ����y�FK����	��Y���ܯ~Zo۝��Ē��X:@cg5l�;o�66"���t��܌r�>�Oe��M��چ��X�v	A�Oܹ��=�Ӓ��C W���8�x��%�Q�N~¢���Zz�}���Lfi��8:8�ͭ��˰�� ���Acĕ�✃U;eZ�g��h���M��xmBډj�\� �;�[��^�W�{Qg.����2	k�,,W���A�J�S��c�䂣)�E�]h3�0���յ���s����zp�W���,#&U�`]L/1Z��ӳN=�����y����Ӌf�}��]b�j1��mN�G�s�cZ�<H��{n/�5a�_	ʗ���#��|�_�?��y��
�\w���E�n�A|�F��4[7�V���V�i�.��9CG��F・��O���+�.�������S��.�������a�q}P�ޚ�wn`���B��C@��A(4�[��}�G�,B٩^�K�(B�E�L��h��:g8z��㣋z�sU'���L�<Bt��5,�5�ե�.���Ӗ#HˎEZ�-HG	���Y��9D�7.*OC���	�*l�y�M�[b��yco{�ٱ�������e�6V`���t�ז2�8o�F���Hn��W�ڝ�7��kW��<��el��W�����Wa�X�m�inKz^��X�'@J���k�R��Ɵ
�v�&���F2���o���[���z��j���*>GqL%���d
:uc}�l�8�^�F�0�����s�q[�O�ϐ��G�͓�i<�	VRh\HT�ӈI�Q�3��:����$���)����y!<`4Ӑ�QCGh����h��T.>����*�L�:���B'J����\�ⳮ[-������$�jl������ץ���5?8 /+�l�����N�^83��t\2.������t�׶+<_�z!~���$�z��#�܋3�) B!�$�rj�݁��P-x!X����Ȍk^6�����Z����JO�w�g�؞��?��?>-����u��pj�O|��.f�ى����������yTv tt�lJv����?j�XOx��H�IC+Oͤ��E7�|���������~m=�K#�~k}��՟z��um����_��>|�x������@ ���t�H1�`�5<�-���)�5G�~YK�.�6����A��^�*Fau�rٯKFXCFM���NC�u}+]//�f�Cw��2l�9�dQ�p��z$�,��X����`񝻇8>?���f��4AVp�;���]�e"-�������!��`�g�-e����Ǡ3_����B����C)���Ȅ@o̴��k^\C��#��:(�.�����wK��{Gv`A�(�)�O�[�2��Cj��lP�6&lA��RҼ*x=�F��K�<S���m�3t��H���R�u�Dz�-�m0��Ȧ� m�����Iy2Y�s��a��y���3x�k�O1��Q�޲C��0���x�s�*jKsIȸ]�y�N%��F� �Η-P9�%���0>�"��e.�~��X�Y"�=ʮ7�|��ږ��R8���VP.�FyU�#�'�8�- ��,@?��B����d��$��8�$,e�Ϫ�C�b��z~��5�(�<���W�������pS��̒s5�n�K^�a5:�G�;vm��kiT�T�`�1�ފ<ʗ���&��[� >�$��\%�����wd&���C"��/��:�+���n^��|a~�<Y}��]��Ve�O{>�X'�u��u4�`�����8�����jx�%8���iD{��<����򦜨+B�M�r}Zn�#�8 n��#�w�������o��P;;X��s�h0`e����k��~�N]g�03�T��z}|p\�>{��M��okG�B�12����=�ש�&�O�;S,"�~����@,����em,OA\�C1p���huQ�'(�=������@�B��h �@�3��E�V��Z�����3�P-#)��[����/�yj�e`:��_�0M�G��	�)�M!F8���u�2�!�ؔ��(썕�>1=�>
/� �pɐ�V����4�	X�m1�_��|��;5D��+`��H���7�f���=�[At��dy��8b�d�
#6)m$����NB�i�7zn�)m����h�P�ܨh`�>o��h�T1Q������]#�W��N����yy�S�<�h6���d������%��sH��F�� � >ǐ��]>d��g\���%b�-W���2��z3�I�'�Y��l;
!ڂ`F��>�!p6%՞��w��I�F��qb$�\5s�"o��^��S��e�К���'�D<�+\��ą&pN��r~���t�-hpl�)_�-ٜ�-
�����W�6
��(����9Z����1�^��9a@~u�xI'��x�ڪm��c��2N�T�G�m���`�hd�tzG�V�3s�Φ=��8$�C�뛈��9[�AYv��Q�3s~�SV�a��Ю��Y�1>�?�塣X���IZ&}BC�ʲ���sߕK��.h;:G��W��h���_`�s0�龨��T}�����?��z}fX����_��[����O�~�Wa ��ـkcG�[�$*����	'�QW$|7��n  ���`\���� <��p�h��>4��Xc��r����^� $��h`~�u�y��׭׷(k�;���$/�
��((�P҇�/2�a^ű)Q!�x����E^[���%`��0�e�C��,t%�٣ȡ��	!wd�҄~�z�� RGۘ��J������'
[�
Z9/^�ӡ�/� f�K�J���|.�d[�pC���R���:�F��t��-c�1^5�����g&̟|f�V.�}�����.�.�l�rs?�!Qo1M�BC�H}�
P%]�l�G��?ޗ[���X���� ��:-N�����i�4R������Z�ѣ��r�Id�T6�b��[�Y?��=�_��(J��+�b���Q�����}6`TG6#6�Pe�Fe�3&��mgKy�R�lFڬs��:9O�A���K�B���|9���ժܦu92[W�Z�� ��A�\E�[:dD�mP	��W�.#'��Y`�A$S��d�43����g����Aâ��!�.l��c�Òw�epi�r_p�4�Y��$��
%#aeP>X/qU>q}jC�GP��R6F�h#թ�4�]�yVx�Aj[�#����H0�!�vZ����y�P�axN���R���7��Z���X �����2���������Am�ۭ��ηn�[sg����@��ژ���7o�N��>�ܮ��^����A*�:s��)����~B�JK߅T�GI���E��c$�`c�5#Wi�K�C oǀ�Ü��퟉t�,���Ͻ*�PB]O�[��4\B�,[���S��wa�<��A��o!����<C��E���xA"�)�(���ZX�_P0�]ŭh��=W��b}�)\wv;;�r_No��#������a��L��9?�c�z�N:�z�ΣGH,oY�{�^����=�ѥpCC8F�FP����J���$p'��"��;m A93�R	�d�U~DC�$��
��R�A*�L��0�e�G�w8�'Q�D�D�.��9�0V��W'�SN�e���[��P$��Wa��변��Dˈ;�G�7#]T��`��rz�yvM>��K��phL�8fY�&xҬ
��A��l���i�s��
WW5��Q4e��p'����$���e� ��m��]�b����E#�:��:}�3?_����Y�E-}��d�$q�p�z���|C�T��-0d���3�iG��Ԅ���h�T��r��m���#��,�'�䬁i�im�O3h?�K?����K,����VnT� ��gI/�����
���Q�[��κp�.�Y]��5ҕ��|��Lr� �ӗF��7|l�k�V];!x>�מ/[3��F���'ڦ�c#��?<���'��O�_�^��:\��?�Z:��������fM�3��� ��,��g4�9���#<4�(P���/�40F@
��R>�ѹq%�XI����c3,�;m���������:�@�J�%�0U���:�c)	b4��my�@%=uX�<k7m��q�>�8G�!~���kHyo��V����t�B5�-us\֣i޳�4�O��ƈF#�mi,^�/m�`��C UJ	�~m��Wgc���[��3'�"��������)08�	d�33:�S
��Q���0��6(���4ki-5�Cw�uHFF9��aL7���|r!G���3L��i�ޣnq���o G��GN�g�`�9ɓ�p%��7�s�"W��|���K�l��rLY������9&;3t�1�$��hWꤜ�'�k�m����t��/���=�����HO��=�9�Ce˩��f�|�HF����� 4>ޗ�/yo[�m}����k�OX2��DЗ��`xL�|�)r�3"ș����j�Sޝ��Q�L8�Hs	J�W�?��	���G]N�Y����W�I���sfs�Kݣ��|�6e��L��`�Q��`�{�)��QL�$J�h���IG ��i��ePj� ��ܺ����)�Q-���ݢ����$�}���J��:cwg��ȇ��3��A��)DT�0���_�_�/�Jm}Ы������E�����a�!֢'4E�0�u����BR��yah�g�Q��(�)7�[ii�ɋ�����{����ΥiL�R�dl��>t�(�N���FT;�ɂ�T�y���#�h��� w,d�咉���N:��Z}��W),�N\O.��L{U �f=�����d(��||>3԰kP�G�D����(��U�x{���o�(F�eXLd��r=��2#őh�!# ����Vk�R�S�T.�W��Ӹ��y�z�6.k�o����v���l�i�qbò�1Li��i?p['�nd \�bQy@R��e��`�a���촖k|7��h�ҏ�پ�G��p��Ӥ��M��>�#�0��>Z�1��|�c�,��T>�E�/$��HR�"�Ȫ��1����$Q�Z[�Q�S�C���z[_M����ƊՄ�(I�[�52ΓD�ͪ���(	����eZ?i��-7ἹЦ�?��	�)e����F^�8]���%>�"Z�%�n�Ȩ���p��9�3��S������W�'����\P,FpC��>o���#n�Nm����-�ёdիpV$i�	L�@OšG�Γ�e�N����:�o�yT!���$�&�F���J	:78;yFNu�BZ	���o&uz��W�8�?��߭��Y�5����>igx>���H�_W�35��!�C��p�ƹW�ھh3���1�F��;`Xf�%5)4�hW�^���Z>��!��Ú��~Mp��s��o�c�-y����E�\.5�ʇ�Π�oR:�tsJC/�G�f.�=5���#�#,�pY��`���8	C���k˛@��,s�������I����g��x�\;tɩ<�@ȥ`�Q�R#�h,^6�V�0|i�~0��K��N/������a����C8���/�fE1(x��؂xe�l�8!8�	��y�Nm�d �
"�2N|�PX�6�8aM�#N�o�w����W�#o�#,�F���n�QY�	�LC����|͑�_������k�8�!����l�)}V�;Kv���Ԏ@��	�V�q��9�:����ht8j��n�@��u�ȉ��b������sx�H�|��>k?��mP	�S�u�Hv�x��x����lun�0q0�Ȓ#�%���B�:���@œ~;g}��6]�g�u��f�(��rh<�&V�k�>���p�MA�@�-�h�b�o2'�
0g�����	u��f8<k+
51���j�$�fF4�(���}c>�t�m�%��He��8�t��sd��ӑ.��Vʧ;��tdE6��2���չ�t�b�'�!uqһ�\a�B��%t�;�qN��� ����Ƕ0��̈3�@e���Xy�?�k���,�{pp�^��y�Kˋ�i�(�E($p���t��.�S��YW�9����xDf)�|f��n9��c>2�	VIY=$o���v�R�s?��9q�錗��e䄶u���v����'���}��z�A��U��Ԋ��}�X�6.u���#>�s��o�$��� �\��D��)�'�~{E�KT�P�,yV ��?���A<T����}~vY[����ZY�c9n���jB�'圮��2#	D|�ѐ�]f��)Z�r߇�SP����*�7^��d�s��{H�B�2A��"04�2U�Qs���'s�0�b���6�m"�n;�h�4E(�� ��R���~!���j���<�N����C:��g�m���p�<�.Xp�k��C.�΃�*-��t5^�ɚ���Hf"e��oEV�������M^b�� #mR� ��h�q����!�����sq��ģ��_�)�>#�H�n�>��(���:��b��w�^��.噁.*���Tʋx5Og�m�>���u�n�(ʳS����Qq�w��b�61�������bX���O�w�f��}� �5�'��un��[(�o^_����(���i���w��"���\�����k���=w
ͣ���Q���T�@�QM�b�ĳ�~`��������{p���e�"��?�.�o�ot�t�v����}��׫�~�N���`ۥƄc�R�C���K=�u⭙���2S;Ǘ��W]���f.�O��Oݾ�RQ��J��7�j��K�꠸O������^B�����|9�sN������f�J���G�{��N�,�\G��v�v�-7��'��׆Jo?32��2�-�P�UD"B>C^?�$s�|N�W?D��s!��J)|p++1���%��|;�!]��fbT�ƩO��~$�|U�9�s�Id[�?�K��m�����e��Q�����<�m���|t�C	���9]��yr�����9�ݹ�<�!���q`y�DY,��@w�V	� �����}���� !��~�p?(�;R����ݤP��4**@�x�jax�x��F�QFJ`*BJC��QG�0�Օ��Q�
ENC'5t��Oe��I'�C�	*^�
|~q>L���QepBg��)��Є���fY����l�
&����Эz܁[���8T�S8���*��31B�#g-x�'Evp���%m�|@��'���RF� $��}&:D^VT`�
!x�3`8��#�����i���Xvm%��zypL��,�ܛ��M?��!t�(����~?�45ajp,�r�FAw,;��g��Ռ_��j�l;3�fz���[��� �E�/��������s���4@	I3��>�#O�X'ڊ�� !0�5�z"���ݐ�����_C+��QX3(�ii=��ٽ���8�5D��y,탊�~���N~�zƍu���*��E����@0��x�nQ%����D��z�R@�a�2e�|*P��Չ������!ݚlIwAH'eT��'�K�l��w�T�jA[�57�(�5�ũ�6����^�2Η��/K�k���¥u�><���z�!|?�/�}1u
Y��B�I��1��{�����e�?�}՝�礱޼��?��6�]����h@?�!y�]`��9���(���E��iC��{�o�����I&Iq�Y0��*����|��v�a=����|g�Bw����vBk�cX��c�Q����a�ҷ�%��]�)��hi���/��K�Z� ��q�wy�
;�:ǶM�X�no��D�\��
U�~��L2�=�b|:��u�o�����{�S���V����;R+��y�U����r�{�$�4$��%;"��l�F�#L���=J&Z2p�E𞻽ڙUN����S�Q�!W �*�Hd�A��͌���VFA���Q�<�\Rp���ü����,ŋhU���Ԣ�F/��e�ӼQ\�����e������6��HpԸ��<��{M*b��@��lxL�j��*�]n��������^da5]��Q9�V(
�\e{���ߊ?����wDG�MMa�4�*Yk�����`�Kq�:�IGH��A�7��V�5܉�A\�U��,!����'O�xd����L��Gً[�'�͔��5G�U;`�5�NI��vA����X/� :�!d[!f����J�7�X��:���9F�%g0Ps(P�|Lۥ}��=FH��m��'e>��gM�[~,��,O��i�<)gy�/r�g�x��S�̣���,�M{�Ӵ��.Y�m&]d+��ڠ���
EZ�A~�xڦ1��ah5����9��TrQ��iT��#��	0�mW� ��8`��`D4��-i�f���t���L���Vۥ�wt����ɏ��T)/��K�w���Vb��֧����]�eQ�k��;��S�e^�B���4 !�:X)!�֨�g����W�Z��.i�B�<�i�z���3�D�!��%9�T��9p�Π%���/ur���֕�Eh����]�S~�F�����:����e��v�X�6�8=u��ޣ�SGzv�!�	��W�e�
[f7�Sà�:�� 
?uI;ꉗ'.�|�L¦�C�ډ$�J�	���C�b1Z������2LnX�^`cft.n��,�l�M�ЎqL1A��D|y�vI���V*�30��.�M"��%t�v
�y��*E����*TҊf��:��գ`�{�C�F�NM6[�JH�8�ь�z.�z1t��t�qܑ�@B��"M,���4�p�b:�x�x�s�����G^�w���o�R�͎H ������QZ�*��Ȝ����͟=��L�M��veB�t,C�*����O�L^�<#K��y�}i���ʉ�8M���W��i���@#G4R��	�drw����r`��]E�M�!=ꏼA^�D,|��&��6�q*����ψ�&��zB'	"�Vakxm���IhLT��� �Qp�{�&*��Y&zۺ������Ƥ�S{�'�uT�!�pi���qor˨��,?��gL8:=��>g��i�H�Ǝ�}qHo���R\�8]��0�3:�� +#A��B�֦�m�:Q��a�K=E�h�vZ�r��8���Q˥�N�xlO�0�%>�Qo+K�mx2�Y���/��HF��ʈ[�{L��3�# �!Od	<�8��^�L�4���H����K����9��4��Lu�o_�O���eC:�̙��C8 D��������a��lp:�%�*�C1����ɈPm�$#d��s� ��i��¢�J��xNR^X�ğ�*=R�$�S�MH�A2�pB@2�0q�Pڭr2BҸ��ad`���I3��ST��q{�IC�����2� ,=?�H� ��4N��a\�_=��y@��l1E��ŨB����b|R^�`�L�I��2+#_"����6ix�o�,����`G��v�Y2�I;ۮP[���k^~����I���0"�7�vq��q�v�GEb�nGp��f�e�H<���#]3��6GF��K�7�`$�-q�QT����G8~�{L��m&��?�\�#�L�|���l�0N1R`|los�4<���.��&�N���%uHX1h��|stb]:3;�J�"<Q�!��#��Eϭ���g�6�,e�:���F>Qr�����k�����IG��Ȇz	?J'tkxI��E�Z2�ȸ�4��i�����Gޤ>��_�q�y��Q:6�9	 	�2�=h�oϬ[�}��@+�u
'6)�	�s�5�l�K�1_��"��E�lG�0zm��奃2�.�S�2��\��Y��ӴS9o2d��䇣۫�p�����xDƅ(�	&&}�<&(�Ӡ�E>UW��z���4;|3=�Jz(?A;A��϶y�О!6\�wN�v�mb!���d�ۯ���D�ᜍ�Dt��Q���vR��*�x�t������ a#Ǟn�^6Ld!�L�aI�C�w�a�D!
��������s�Pّ�gCi���x'�M;��<mA�X8��}�������yN���im�,�ܦt�+|a����2֯75���s:�^Zc��1�����v�q�<�j{���	�v��%��p�&G�����Zû�<Q 6|tm�PK�i����>��e1>
T�H��q��1��2J��JxyMq��N�|��ҕ5�9���4=ϴ"�kC�8�������s��m�#��_�K�VF�k;U��F[�aj��
�4#:�r�|�Ea�딗Fd�RGdzg����q]!����:Ubv���:������H=��*��i@�n��ӌ[3
_�\�Nڥ�RN[n��m���M�4m7a:%;6y6�4%a��g��4ᇀ��i�e\�4�A�J>�Xʯp��u
#��g��~볶�ɮ��(Vdέj��ǈg�O�4�#K�&� �c�����ayy�������H��'�?|��`kl�͖��6���O�R<�����q�x��,O�K�U�d��8�y�3Z��-�Os*��?��u�t������s���N�x�3v�ѥ�+�Gp�څT��#��㠌)�i Z[�C;�CQ�#��N�>�᫴���Q�B%����*H����|Rwn��v,�X<U�;G�W��t���AS�0e��0�d�����ݼ�b^N-)�1>
�xMe�M���9e���+C;�J���'L�ɒ(��O,m�2�<L�S IB8��9ZQpQp>�Sѓ�:T��2�+t�gk�M�c��AFJNC4�hY^�Tp�$�8;�dE�a��n}�)�f���/q�J��X�SE#m�,�hs��|��d�W*�8#Û|�'0�!��9�y�^�'���q1��1� u�7< t1����Ҷu�I>��[p���&uX�iN覲톣��5D)PW�(��+��j�^�V�r?r+�(i�H�s;E3����6C�K�sߞ'�+�^U�s�PYk/iҤ9C��/ب��@�㸉�x��E�"�#�I#ZS�]�C{�:�
M�V��Od�h=FZ�";�	��k��1eGii8������y����ǫ#]�� �f݉9���<6��I<ϣ���"��8B8~�uXW���&�s�3���87\�e����^�*~҇v�,���^#:�M҈[z�ʄ#�о5:r��e�}�{��e�{�3e�V�eŪu�+���f(I��M>|�a��m���$R��w!�F��s-��qZ��2=���@C��/�G�1_��)�	�)��O=��6���L�>~�ҍ)mg��^��S:B�  ?�j!@#�^I�?=5a9����Va�he�!hj�,K��� |<��BT!D	ڨ���r�1Kd9��{Yl1m>e#l�Nl��?s� %�}�>����F��0�u��7�XfJ�Q��L� l�|����y�t�LsD/�yW�z4�
��H�7ϼl#���FY�5B��֪$,�I]�|���Z���h^{�K���M�g�8Q�w(|WJ����GICo�{>�g�S��ɔt��_<5�cYS�5@�Q�/˙?�R�	�vn0ke��3G`���ШތZT��(_y���+L'��d!��&�A堓�3Aq�����im�M򋟰�e��oNR�g�r���Z�!�����x��Z�=��
д�w9����1ā�4�2���&
G�m�Ѿ��2y��i��~�o�:�)�9�v+g^o��q��y��A��"�ߜ�pE�8O����7��>�Q��%��	~=�&m43v �cC�(]��	:yo0�'פ��Q��~0���Ȟ�^q5-#8�S��i���n�!�_�����4�}�8�ԗ~�_�1���y��Y�r��58pO�c�p#%l���~ϭ�6�؀\�*Cd��'M�i�ԁ���?X�LIEc�SdXg2��d7F�:����pu	��\��~��@l
�|�[H*`��?#fX3UDt��F>ײ����%M�!��φ��V��T��)cǇ��XQd��i�U��)����h#��9�5EJ�"o���1b�E踥�� ~~Z����b��xY�Y�h��S�� (���
m� ��:f�z�>Rbq�"�
mo)�3�Te��E��,W��8!�\���$��<�K�n�L9σB:P~����vy�B��H5XЙ���2℀Ű�k��8�s�G
4.�C3p��[��y��#�N���^Ey���O�m����6�)/!����j:@�L=�V�Bx�NFeĕ����"�*���3�?NP��i��� ��P�rM>a����)�Y��^.s`9E��sRi�!*���Z����t��L����G���͋���M�A�2���un���o�I�ȍ�N��Pd��a��S�9��>�:���`@7i/��گq�@�.i�m���!���6zo�*�B���h�G�s��m�Y����� ����(�\G޹��6���GDC|�iF�\�h��)�]�f��j�Ƒ8��<�p�h򓦳*��w�{�|5��E��6�ԭ�rK����AjӍ1(����� ���8���yc���K�@#����!����bxB=���/^��f1i���c�gj�'�]�'<i�rK��%�+��6�/��x���H)����VSh�Ul�ͧ�9wa��b�$P���i�>z=?��� /��ڡ4�<_�!AZ$9��0F�4/�ՇwQ���Y����R�#���%<��o�������P蚒�q�K�
��� �^'m�}�t)�0���$*��檿��#��|{�;�����ySc���H{�V����z�~)�2r�u(1ĴS����Ŵ��� �%��/=B��4��i/��G���QD���+�=�/�#ժ�~��G��6鏤潑�vi�͛|��.���j�>逪J��$q�F��/Q��N�#���R��V6�@���F�xR:��S�V��lt��	2^#_�[�����ʷ<j�]���#0#g�����x�����74Ά6"����_C�Q�}:�Qd��zLp�g+�-&�ڗY�#��U�#�l�t�*�3e�G�FVF����6�&�J�%-Z��&��K�'��H��O��υ�/�����M�<SJ�%Mކ�<c��h(��s�ݥ16�~Ã8��΃�QSǵ�U�.�f�gb'T�r��<IQ���mC��t͸�c�Ae�d���X���m���נ�����'bs$�Y+�yJea�4%��/�䧼���´MvE�cF���6�w�t%����M�ͣ4�i�rԧ�R��?���&������@9�    IEND�B`�PK   �cU!�`�-  �     jsons/user_defined.json��]o�0��J��`��8wQ"U�֮k�i�MĘ�Zj��UQ��>�4�6�Ԩ�
���x^X�fU0mm���֙��O�k[�0� �8���+����zq�=uk�?�P���<�~
��@�����#`�P&1�(pRPM��H��dQ(#R���U�t�엎ߚ�{�L����]c��n�����=�u�uW�(�x\�4�u��V�rn(�!C�a�|�0��r�v�ݓh��ц�U~�x��uem�F��2����2�%��8���a��F���t���S�����J/�e���fvO�x1?C'�GgC�@�o���N�g�*�0�����n%�ӥ�F���r_���ȝ�<G\���H��,�t8CY�)2�q�� w>BnEJ�q�)�(b��+��b�I��$B���7�������~��������b8�\@Y.��8��5ƹlx��=��]����g���1�Zb�H�`�݊�DQT$k�n0foIT>"Q$|�xz<R��(�	�T <�\@�$a���mꀧ�����W|9�c���	BP D�~HC]�~����PK   �cU9_���P  �[            ��    cirkitFile.jsonPK   �cUs�7+5J  dK  /           ��Q  images/6c71542d-16cb-4630-930f-71c4de5e1144.pngPK   �cU����:  ;  /           ����  images/71057ff1-f3c2-49c6-8a17-bf9e68e09ed9.pngPK   �cU��g� s� /           ��g�  images/d4dd056e-e2cb-4614-accb-0aa130e74534.pngPK   �cU!�`�-  �             ���t jsons/user_defined.jsonPK      �  $w   